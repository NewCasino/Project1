﻿ABN AMRO Bank
