Det nya lösenordet får inte vara samma som något av dina tidigare lösenord.