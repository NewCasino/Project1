﻿Formatet i fältet är ogiltigt. ( e.g. FI2112345600000785 )
