﻿Upprepa lösenord här
