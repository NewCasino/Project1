﻿Laddar
