Uttag av pengar direkt till ditt PRZELEWY-konto