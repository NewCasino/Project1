﻿Belopp att överföra


