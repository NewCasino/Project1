Summa är utanför de tillåtna gränserna