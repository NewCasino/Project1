Stäng den här dialogen