[Metadata:value(/Metadata/Settings.Operator_DisplayName)] – Ditt användarnamn är här