Kredit kort