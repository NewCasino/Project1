﻿Tårtpokerbonus
