Lördag