﻿Inloggning
