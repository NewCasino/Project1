﻿[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Meddelande om ändrad e-postadress