Giltigt från