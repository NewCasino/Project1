Uttag av pengar direkt till ditt VISA Electron-kort.