﻿Mobil