Gäller fr.o.m. : {0}