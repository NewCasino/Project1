Region / landskap