﻿Sport Vinnare
