﻿PayU