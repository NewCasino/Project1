﻿i-BANQ användar-MID lösenord krävs
