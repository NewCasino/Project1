Du har uppdaterat din profil.