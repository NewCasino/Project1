En 30-dagars självuteslutningsperiod