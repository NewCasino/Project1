Voucher-numret krävs.