﻿Är du säker på att du vill avsluta denna kod?
