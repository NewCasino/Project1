﻿<p>CEPBank:</p>
<p>När pengarna har mottagits och klarerats, kommer vi att kreditera ditt spelkonto. Du behöver följande uppgifter när du gör en banköverföring till ditt spelkonto.</p>

<p>Gör insättningen till
 <ul>
 <li> <strong>Kontoinnehavare</strong> : OddsMatrix Ltd</li>
 <li> <strong>Innehavarens adress</strong> : Vincenti Buildings, Suite 713, 14/19 Strait Street, Valletta, VLT 1432, Malta</li>
 <li> <strong>Bank na</strong> : Bank of Valletta</li>
 <li> <strong>Bankens adress</strong> : 86, South Street, Valletta VLT 1105-Malta</li>
 <li> <strong>SWIFT</strong> : VALLMTMT</li>
 </ul>
</p>

 
<p>
Nedan visas IBAN-numren för vardera valuta
<ul>
<li> <strong>EUR</strong> MT25VALL22013000000040018502408</li>

<li> <strong>SEK</strong> MT11VALL22013000000040018502466</li>

<li> <strong>DKK</strong> MT34VALL22013000000040018502440</li>

<li> <strong>USD</strong> MT04VALL22013000000040018502495</li>

<li> <strong>GBP</strong> MT73VALL22013000000040018510759</li>

<li> <strong>NOK</strong> MT73VALL22013000000040018502453</li>

<li> <strong>PLN</strong> MT73VALL22013000000040019112062</li>

<li> <strong>CZK</strong> MT13VALL22013000000040019112075</li>
</ul>
</p>

<p>Observera att vi inte debiterar dig för insättningar via banköverföring men vi rekommenderar att du kontrollerar med din bank om eventuella tillkommande avgifter, intermediära bankavgifter, som kan förekomma. 
</p>