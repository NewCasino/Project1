﻿{0} tillgänglig