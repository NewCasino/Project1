TC Nummer