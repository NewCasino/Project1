﻿Inloggning med användarnamn är inte tillåten för verifierade konton. Vänligen logga in med ditt NemID.

