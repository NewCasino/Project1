Med ditt Visa Electron-kort kan du snabbt sätta in pengar på ditt spelkonto via Skrill. Du behöver bara registrera ditt kort på Skrills gateway och så snart ditt kreditkort har verifierats kommer pengarna att föras över till ditt spelkonto, säkert och omedelbart.