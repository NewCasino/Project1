﻿Master Card