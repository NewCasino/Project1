Jag har läst reglerna och villkoren