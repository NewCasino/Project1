Ons