Begäran om allmän support