﻿Ladda Saldon
