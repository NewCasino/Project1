<em> Detta e-postmeddelande skickas av kunden på "Kontakta oss" sidan. <br /> Svara INTE på detta mail direkt! Du hittar kunden emails nedan </em> <hr/> <ul> <li> <strong> kunden E </strong>:. $EMAIL$ </li> <li> <strong> Kundens namn </strong >: $NAME$ </li> <li> <strong> Ämne </strong>: $NAME$ </li> <li> <strong> användar-ID </strong>: $USERID$ </li> <li > <strong> Användarnamn </strong>: $username$ </li> </ul> <hr/> <pre> $ INNEHÅLL $ </pre>