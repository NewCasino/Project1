﻿Jag har läst och godkänner informationen jag har fått
