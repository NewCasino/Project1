﻿/game/gamerules.jsp?game=roulettemini&lang=sv