Ditt personliga ID har redan registrerats