﻿Pott
