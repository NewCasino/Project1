Otillräckliga medel.