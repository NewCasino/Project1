﻿/game/gamerules.jsp?game=sevengoldscratch&lang=sv