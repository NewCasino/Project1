Visa alla