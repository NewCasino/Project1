Ditt konto ID måste vara minst 12 tecken