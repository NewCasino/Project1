Address rad 1