Ange din e-postadress