Visa dina favoritspel