Kontouppgifter