﻿Vänlgen välj ett kort.
