Är du redan en EntroPay-användare?