Välkommen {0}