﻿Vouchernummer
