Den här transaktionen har rullats tillbaka.