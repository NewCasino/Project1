Spela {0} nu!