Lösenordet upprepades inte korrekt