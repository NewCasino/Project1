﻿/game/gamerules.jsp?game=eldorado&lang=sv