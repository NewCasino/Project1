Lokal banköverföring {0} {1}, internationall banköverföring {2} {3}