﻿/Metadata/Villkor
