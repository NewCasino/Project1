Gör ett uttag direkt till ditt Moneta konto