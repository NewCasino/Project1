Du spelar i underhållningsläge.