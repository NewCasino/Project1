﻿Deltagare
