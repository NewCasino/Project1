﻿Avbryten