﻿Cake Poker Turneringar
