﻿Välkommen
