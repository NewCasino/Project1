Välj ett konto