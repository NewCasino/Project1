﻿Ditt uttag kommer att behandlas så fort som möjligt.
