﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)]: Prisänkingsmeddelande
