Gör ett uttag direkt till ditt TLNakit konto