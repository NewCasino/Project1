Innehåll