Lösenordet har inte upprepats