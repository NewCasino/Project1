Personligt ID-nummer