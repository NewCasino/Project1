Insatsgräns