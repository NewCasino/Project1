﻿Vänligen ange ditt Konto ID.
