Gå till vår Sports Book nu!