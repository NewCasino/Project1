du måste logga in först, innan du kan spela med riktiga pengar!