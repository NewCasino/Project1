﻿Observera! Vänligen skriv ner den genererade tillfälliga koden som presenteras ovan, (Gilltighetstiden av koden är 12 timmar)
