Lägg till pengar