Gräns: