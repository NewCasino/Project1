Du får inte ändra e-mail på grund av ofullständing profil. Du kommer att bli omredigerad till profilsidan om 5 sekunder, var vänlig färdigställ din profil innan insättning.