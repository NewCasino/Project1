﻿Land Blockerad

