﻿<img src="//cdn.everymatrix.com/Shared/_files/Meddelande/skickat_mail_24x24.png" alt="Skickat från mig" />
