﻿UK Gambling Commission Villkor och bestämmelser