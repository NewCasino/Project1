Du måste logga in för att rulla tillbaka uttag.