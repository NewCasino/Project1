﻿Land
