﻿Klas Poker Bonus
