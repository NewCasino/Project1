Tack, din begäran kommer att behandlas så snart som möjligt.