Min favoritbetting?