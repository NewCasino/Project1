﻿Skicka ny verifieringskod ({0} seconds)

