﻿/game/gamerules.jsp?game=lrroulette2french&lang=sv