﻿Check nummer