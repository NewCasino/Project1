Kontrollera att valutan och beloppet ovan överensstämmer med valutan och beloppet på din IPS-voucher.