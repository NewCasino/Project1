Bank/kredit kort