﻿Casino FPP