Gör ett uttag direkt till ditt AGMO konto