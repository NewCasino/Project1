﻿Vänligen skriv in IBAN
