﻿Tillgängliga turneringar
