﻿Jackpot i 53