﻿Lösenordet måste innehålla bokstäver och nummer.
