﻿videokolikkopelit
