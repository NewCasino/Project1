﻿/game/gamerules.jsp?game=maxwin&lang=sv