Självuteslutning