Uttag direkt till ditt MONETA konto