﻿Kundtjänst
