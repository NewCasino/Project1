﻿Hem
