﻿<!—Infoga logga här --> 
