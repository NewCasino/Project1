﻿jattipottipelit

