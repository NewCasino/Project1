﻿/game/gamerules.jsp?game=lrblackjackflash&lang=sv