﻿Om Nordic777



