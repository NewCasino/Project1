﻿Alla Överföringar
