Gränsen har tagits bort men den gäller fortfarande fram till utgångsdatumet.