Gränser: