﻿Omaha