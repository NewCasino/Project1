﻿Fullbodad
