﻿Vänligen skriv in din väns användarnamn
