﻿Alla Amerikanska I
