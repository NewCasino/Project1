Efternamn