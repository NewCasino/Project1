Låt mig aldrig logga in igen