﻿http://stats.egtmgs.com/jackpot_ExclusiveClub_EUR.json
