﻿Misslyckad