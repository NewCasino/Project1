Mottagarens telefonnummer