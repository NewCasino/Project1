﻿Deposit with Bank Wire