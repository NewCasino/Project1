Läs villkoren här