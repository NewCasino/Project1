Registrera ditt konto