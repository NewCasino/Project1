Ämne: