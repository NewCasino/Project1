Betala per telefon (Australien)