Uttag direkt till ditt Poli konto