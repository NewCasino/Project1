Antal vinnare: