﻿/game/gamerules.jsp?game=luckyeightlove&lang=sv