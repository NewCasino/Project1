﻿Vänligen skriv in clearingsnumret
