Betala per telefon (Nederländerna)