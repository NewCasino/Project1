Uttag av pengar direkt till ditt VISA-kort.