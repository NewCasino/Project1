﻿/game/gamerules.jsp?game=jackhammer&lang=sv