Ange ett giltigt datum.