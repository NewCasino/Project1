﻿Spelpengar (av Dotpay)