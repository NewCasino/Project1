﻿Steg 1. Logga in manuellt på <a style="text-decoration: underline;" href="{0}" target="_blank">din onlinebank</a>
