Uttag direkt till ditt Clickandbuy konto