Du dirigeras om till giftcardempire.com när du klickar på Fortsätt