<p>Kära $USERNAME$, <br /><br />Tack för att du kontaktar [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br />Detta e-postmeddelande är för att bekräfta att du har ändrat din personliga insättningsgräns från $LIMITAMOUNT$ $LIMITPERIOD$ till $NEWLIMITAMOUNT$ $NEWLIMITPERIOD$. Den nya gränsen kommer att aktiveras på $LIMITEXPIRYDATE$. <br /><br />Tveka inte att kontakta oss om ni har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p><br />Kind Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kund Support Teamet</p>