﻿[Metadata:value(/Metadata/GammingAccount/IGT.Display_Name)] Kredit & Debet

