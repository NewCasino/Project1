Summa kan inte vara tomt