Se föregående spelsida