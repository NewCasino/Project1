﻿Ta det!
