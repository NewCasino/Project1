Från