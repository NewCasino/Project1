Överföring av pengar direkt till ditt EcoCard-kort