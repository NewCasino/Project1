Välj sorteringssätt: