<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Syfted med detta e-mail är att bekräfta din personliga förlustgräns $LIMITAMOUNT$ $LIMITPERIOD$ kommer att försvinna den $LIMITEXPIRYDATE$. <br /><br /> Var vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p><br /> Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>