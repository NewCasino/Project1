Uttag av pengar direkt till ditt Neteller-konto