﻿Ange lösenord här
