Din överföring av pengar lyckades.