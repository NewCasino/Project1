﻿jattipottipelit
