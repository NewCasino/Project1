Jag har en bonuskod