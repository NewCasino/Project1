Lägg till ett nytt spel