﻿muut-pelit
