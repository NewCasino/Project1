Vänligen välj en säkerhetsfråga