﻿Vänligen ange ditt mobilnummer
