﻿Filialkod