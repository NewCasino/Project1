Direkt e-banking