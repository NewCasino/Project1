Giropay är en online betalningsmetod som fokuserar på den tyska marknaden.