﻿Beskrivning
