Uttag av pengar direkt till ditt GiroPay-konto