﻿United States