Välj kompis för överföring