Rulla tillbaka