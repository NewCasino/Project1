﻿/game/gamerules.jsp?game=wildwitches&lang=sv