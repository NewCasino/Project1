﻿Vouchernummer måste bestå av 16 siffror
