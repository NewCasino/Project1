Neteller Konto ID