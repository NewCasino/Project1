Uttag av pengar direkt till ditt Georgian Card.