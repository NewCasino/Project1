﻿Minimal poäng att hämta:
