﻿Kolla vilket fantastiskt utbud av fotbolls-, basket-, handbolls-, tennis- och ishockey-matcher vi har i vår Sport-sektion idag! Vi har de flesta av världens sporter och tävlingar även utan live odds.