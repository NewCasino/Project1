﻿[metadata:value(/Deposit/_Index_aspx.Button_Confirm)]
