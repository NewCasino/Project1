Kontoutdrag