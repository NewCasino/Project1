﻿Jag har läst och godkänner reglerna ovan
