Ditt svar