﻿Saint Kitts And Nevis