Välj en säkerhetsfråga