﻿UIPAS Konto ID
