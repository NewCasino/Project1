﻿/game/gamerules.jsp?game=retro-funky70&lang=sv