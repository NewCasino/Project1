Överföring av pengar direkt till ditt Intercash-kort