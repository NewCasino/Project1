Ändra...