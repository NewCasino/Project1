﻿Insats
