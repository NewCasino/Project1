﻿Överföring

