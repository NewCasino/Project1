Romänien, New Leu