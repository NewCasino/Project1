﻿scratch-cards
