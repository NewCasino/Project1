Välj ett betalkort.