E-postadressen inte tillåten