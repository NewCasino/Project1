Utfärda ett IPS-tecken och för över pengar till den nya vouchern.