Du får inte göra en överföring.