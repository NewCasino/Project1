Dealerns kön: