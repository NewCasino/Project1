﻿Referensekod
