﻿Kasino Hold'em
