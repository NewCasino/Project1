Du har avbrutit transaktionen.