Ditt lösenord måste bestå av minst 8 tecken