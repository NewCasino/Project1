﻿/game/gamerules.jsp?game=bingo&lang=sv