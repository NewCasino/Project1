﻿Sida:
