Detta fält är ogilltigt