﻿SinglePlayerPoker