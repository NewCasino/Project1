Insättningsgräns