﻿Neteller(Mexico)