﻿Avslutad av ATM
