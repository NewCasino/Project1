﻿Singel Deck Blackjack Serier

