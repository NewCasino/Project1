Referensnumret