Vänligen fyll i mottagarens turkiska National ID