﻿Visa endast {0} spel