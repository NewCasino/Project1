Inledande vadslagningskrav