Det här fältet är ogiltigt