﻿Insättningsgräns
