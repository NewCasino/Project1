Aldrig