Välj ett konto.