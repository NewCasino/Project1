﻿/game/gamerules.jsp?game=piggyriches&lang=sv