användare