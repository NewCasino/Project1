Vänligen ange medborgar ID