Vänligen fyll i bonuskoden.