Uttag av pengar direkt till ditt Baloto-konto