Direkt