﻿Inställningar
