﻿Valideringskoden måste bestå av 6 siffror
