﻿Dubbel Exposure Blackjack Serier
