Gratis