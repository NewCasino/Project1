Vänligen ange din adress