﻿Välj ett konto
