Öppna spel i helskärmsläge