Ändra