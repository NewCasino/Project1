﻿/game/gamerules.jsp?game=egyptianheroes&lang=sv