Belopp som ska tas ut från {0} konto.