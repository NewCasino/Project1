Vänligen ange ditt postnummer