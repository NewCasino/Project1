Till en kompis konto.