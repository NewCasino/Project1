﻿NYXGaming