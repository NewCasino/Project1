﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)], Självexkluderingen har avslutats
