﻿Tack, din förfrågan behandlas så snart som möjligt.
