﻿<p>Hej $FIRSTNAME$,</p>
<p>Det här automatiska e-postmeddelandet är ett kvitto på din insättning som har behandlats på uppdrag av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] av OddsMatrix Ltd, betalningshandläggare för [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] webbsida, kommer du att se EveryMatrix på ditt kort- eller bankkontoutdrag. Dina transaktionsdetaljer visas nedan.</p>
<ul>
<li><strong>Transaction ID</strong>:$TRANSACTION_ID$</li>
<li><strong>Date time</strong>:$TRANSACTION_TIME$</li>
<li><strong>Webbsida</strong>: $TRANSACTION_SITE$ </li>
<li><strong>Kvitto</strong>: utskriftsversionen av kvittot i bilaga.</li>
</ul>
<p>Har du frågor angående den här insättningen, kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a> hänvisa till transaktions-ID-numret.</p>
<p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet</p>
<p>$SCREENSHOT$</p>