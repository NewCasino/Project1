﻿Duplicated vendor limit rule