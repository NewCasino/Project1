﻿Deuces Wild Video Poker Serier
