﻿Hem Bonus
