﻿/game/gamerules.jsp?game=hrhilo2-3c&lang=sv