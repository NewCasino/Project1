Beloppet överstiger gränsen.