﻿Vänligen skriv in kontonumret
