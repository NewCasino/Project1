﻿videopokerit
