Laddar