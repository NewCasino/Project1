Belopp som ska överföras