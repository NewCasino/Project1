﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Ditt uttag har nekats

