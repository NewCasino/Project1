Uttag direkt till ditt WebMoney konto