Vänligen fyll i innehållet. 