﻿Om
