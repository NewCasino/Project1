Gränserna är borttagna, men de gäller tills slutdatumet