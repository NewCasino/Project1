﻿/game/gamerules.jsp?game=hrbaccarat2&lang=sv