Fel