ingen tillgänglig bank