﻿Hem

