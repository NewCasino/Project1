Villkor & bestämmelser