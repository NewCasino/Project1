Nyligen använda kort