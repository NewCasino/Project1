Du kan begära uttag med följande metoderna som finns tillgängliga för dig