﻿Table Games

