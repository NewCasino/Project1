﻿Du måste logga in för att se dina tillgängliga bonusar.