﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Aktivera ditt konto