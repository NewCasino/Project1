Du har lyckats med insättning.