﻿Välj din bank
