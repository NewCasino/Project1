Ange bonuskod.