﻿Bankuttag med Trustly
