﻿Du kan snabbt sätta in pengar med ditt VISA-kort till ditt spelkonto. Ange kortuppgifter och så fort din betalning har godkänts av din bank, krediteras ditt spelkonto.
