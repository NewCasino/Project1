﻿* <em>Bonus på din insättning: {0} {1:N2}</em>