Misslyckades!