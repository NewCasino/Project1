Lägsta insättningsbelopp