Ogiltigt Ukash värde