﻿/game/gamerules.jsp?game=lroasispoker&lang=sv