Logga in