Ditt valda användarnamn finns redan registrerat, var vänlig och välj ett nytt.