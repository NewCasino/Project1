lyckades