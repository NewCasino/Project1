Betala per telefon (Frankrike)