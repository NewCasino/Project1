Dina sammanlagda uttag överstiger 2 300 EUR och vi är tvungna enligt lag att verifiera ditt konto innan vi kan behandla ditt uttag. Skicka följande dokument med e-post till <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>
<p>a) bevisning av adress, t.ex. en räkning eller ett kontoutdrag </p>
<p>b) en kopia på nationellt ID-kort eller pass</p>
<p>c) en kopia på kortet som användes vid insättningen</p>