﻿<ol>

 <li> <strong>Hur gör jag ett uttag från på mitt webbkonto?</strong>
 <p>
Du kan begära ett uttag när som&nbsp; helst&nbsp; så länge du uppfyller alla krav och har&nbsp; auktoriserats för uttag i vårt system. Du kan också göra så många uttag du vill men på grund av lagstiftning mot penningtvätt och bedrägerier som gäller här [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kan vi inte medge uttag från ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]&nbsp; konto förrän 24 timmar efter det att du gjort en insättning. &nbsp; Ett uttag måste uppgå till minst 10 Euro.
 </p>
 </li>

 <li> <strong>Finns det någon gräns för hur mycket jag kan ta ut?</strong>
 <p>
Ett uttag måste uppgå till minst €10.00 eller motsvarande i din valuta. Ett uttag får uppgå till max €5000 per dag eller motsvarande i din valuta.
 </p>
 </li>

 <li>
 <strong>Kan jag ångra en uttagsbegäran?</strong>
 <p>
 Du måste kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kundtjänst och om&nbsp; uttaget inte har behandlats kan det stoppas.
 </p>
 </li>

 <li>
 <Kan jag få mina vinster betalade tillbaka till mitt kredit-/bankkort?</strong>
 <p>
Ja, det kan du, så länge det är samma kort som du använde för att göra den ursprungliga insättningen och om kortet kan&nbsp;  ta acceptera en&nbsp; återinsättning.
 </p>
 </li>

 <li>
 <strong>Jag använde mitt kredit-/betalkort vid insättningen, kan jag begära en utbetalning på något annat sätt?</strong> 
 <p>
Ja, det kan du men vi kan behöva fullständig dokumentation från dig och uppgifter om ditt nya sätt.
 </p>
 </li>

 <li>
 <strong>Varför kan jag inte välja på vilket sätt jag vill ha utbetalningen?</strong>
 <p>
 Det beror på lagstiftningen mot penningtvätt som vi följer och för din och vår säkerhet i alla ekonomiska transaktioner, så utan auktorisation måste alla insättningar gå tillbaka till samma metod som användes vid insättningen.
 </p>
 </li>

 <li>
 <strong>Har ni särskilda avgifter för uttag?&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;</strong> 
 <p>
 Uttagsavgiften varierar beroende på vilket uttagssätt du väljer. Vänligen Klicka här '
 <a href="/depos>Betalningsmetoder</a>
 " för information om avgifter och tänk på att din bank kan debitera dig en avgift för sina tjänster.
 </p>
 </li>

 <li>
 <strong>Hur lång är handläggningstiden för?</strong>
 <p>
 Detta kan variera beroende på vilket uttagssätt du väljer. Vänligen klicka här '
 <a href="/depo>Betalningsmetoder</a>
 ' to see all of the withdrawal methods available to you and their processing times.
 </p>
 </li>

 <li>
 <strong>
 Why is it that a withdrawal to my card takes days while a deposit is immediate?
 </strong>
 <p>
 Vi gör ett antal kontroller och utredningar innan några uttag lämnar  [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] och detta fördröjer uttagen med cirka 12 timmar. Dessa kontroller är en del av våra löpande åtgärder för att säkerställa säkerheten för våra kunders pengar. Alla andra fördröjningar beror på restriktioner som påtvingas av betalningsleverantörerna.
 </p>
 </li>

 <li>
 <strong>
 Vad händer om kortet som jag gör uttaget till har gått ut eller dragits tillbaka?
 </strong>
 <p>
 Du måste meddela oss om alla ändringar i&nbsp;  kortet och lämna in bevis på utgångsdatum eller orsak till ändringen.&nbsp; Ett nytt kort måste registreras hos oss och på ditt  [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto.
 </p>
 </li>

 <li>
 <strong>
 Kan jag göra ett uttag från mitt konto och få dem skickade till någon annans konto?
 </strong>
 <p>
 Nej, det anses som en tredje parts-transaktion och är under inga omständigheter tillåten.
 </p>
 </li>

 <li>
 <strong>
 Vilken uttagspolicy har [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayNa)]?
 </strong>
 <p>
 Ditt konto måste vara aktiverat och ha minimibeloppet som krävs för att göra ett uttag. Vissa restriktioner kan gälla för spelare som deltar i [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kampanjer.
 </p>
 </li>

</ol>

<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Print</span>
 </span>
 </span>
 </span>
 </button>
</p>