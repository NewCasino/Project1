﻿Registreringstid
