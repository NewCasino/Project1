﻿/game/gamerules.jsp?game=knockout&lang=sv