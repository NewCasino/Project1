﻿Avslutad
