﻿Ortfältet får inte lämnas tomt
