Användar-ID