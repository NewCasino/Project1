﻿Välj en vän att överföra till.
