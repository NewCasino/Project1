Registrera