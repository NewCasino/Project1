﻿Transaktionen kan inte stödjas för tillfället.
