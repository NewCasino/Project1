﻿Aktiverar registreringen med användarnamn och lösenord
