﻿ASN Bank
