﻿{0} secunder

