Vänligen fyll i referensnumret.