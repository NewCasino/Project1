Ange Ukash-värde