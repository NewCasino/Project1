Ryssland, Rubles