Belopp som ska överföras till {0}