﻿/game/gamerules.jsp?game=oasispoker&lang=sv