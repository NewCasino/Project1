﻿Vänligen klicka i checkboxen
