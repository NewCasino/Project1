Belopp