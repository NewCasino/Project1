﻿CASHU