﻿Voucher