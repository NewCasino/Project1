﻿Avgift
