Namn på ditt konto