Ändra e-mail