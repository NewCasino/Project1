﻿/Kasino/Info/SpelRTP
