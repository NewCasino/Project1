IPS-tecken