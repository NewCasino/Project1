För att debiteras från {0}