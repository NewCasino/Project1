﻿/game/gamerules.jsp?game=eldorado_sw&lang=sv