﻿QIWI

