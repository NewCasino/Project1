Debitering misslyckades