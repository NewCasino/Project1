﻿/game/gamerules.jsp?game=hroasispoker&lang=sv