﻿Deposition →
