﻿Utloggad
