﻿/game/gamerules.jsp?game=minispellmini&lang=sv