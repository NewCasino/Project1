Visa turkiska bord