﻿Euteller är direkttjänst för internetbanköverföringar från Finland
