Ogiltig säkerhetskod