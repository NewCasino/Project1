Ingen gräns