﻿Clearingsnummer
