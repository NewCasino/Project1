﻿Ditt uttag kommer att skickas i EUR pågrund av spel regleringen i Norge, notera att beloppet kan vara något mindre på grund av valutakonvertering.
