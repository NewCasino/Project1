﻿Överföring ID
