Akbank är en turkiskt baserad bank