Välj din region