<strong>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] AVSLUTA ANVÄNDARAVTALET</strong><br/><br/>VÄNLIGEN LÄS FÖLJANDE NOGA. VI REKOMMENDERAR DIG ATT SKRIVA UT DESSA VILLKOR OCH BEHÅLLA DEM TILLSAMMANS MED ALLA BEKRÄFTELSE E-MAIL, YTTERLIGARE VILLKOR, TRANSAKTIONER, SPELREGLER OCH BETALNINGSMETODER DÅ DE RELATERAR TILL DIN ANVÄNDNING AV SIDAN. VI SPARAR INTE VARJE INDIVIDUELLT KONTRAKT MED VÅRA ANVÄNDARE VAR DÄRFÖR VÄNLIG OCH SKRIV UT DEM FÖR ATT SPARAS. DESSA VILLKOR KAN ÄNDRAS UTAN FÖRVARNING.<br/>ANMÄLNINGAR AV DESSA VILLKOR UTGÖR TILLVERKLIGEN AV ETT ERBJUDANDE. GENOM ATT REGISTRERA TILL ANVÄNDNINGEN AV DESSA TJÄNSTER SOM OMFATTAS AV DETTA AVTAL, FÖRSÄKRAR DU ATT DU ÄR 18 ÅR GAMMAL OCH DU SAMTYCKER ATT FÖLJA FÖLJANDE VILLKOR. OM DU INTE VILL ACCEPTERA DE FÖLJANDE VILLKOREN, SÅ KOMMER DU INTE REGISTRERAS OCH ÖPPNA ETT KONTO OCH DU KOMMER INTE FÅ TILLGÅNG TILL MJUKVARAN OCH SPELTJÄNSTERNA SOM ERBJUDS I SAMBAND MED DEM.<br/><br/>Det här avslutar användaravtalet (“Avtalet”) är ett juridiskt bindande avtal mellan Dig (”Dig”) och [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], som drivs av EveryMatrix N.V. , ett bolag bildat i Curacao, och företagets dotterbolag, efterträdare och övertagare (kollektivt hänvisade till häri som"[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]"). Mjukvaran ("Mjukvaran") och speltjänsterna ("Speltjänster") tillhandahålls till Dig av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] på en ”BEFINTLIGT SKICK” grund, för Din personliga användning, endast. Pokerapplikation och mjukvarand som används på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] hemsidan drivs av EveryMatrix NV, ett bolag bildat i Curacao, som har en Curacao spellicens No. 8048/JAZ i november 1996 No. 41.<br/>Vänligen notera att mjukvaran och Speltjänsterna INTE ÄR FÖR BRUK AV PERSONER UNDER 18 ÅRS ÅLDER. Ingen under 18 års ålder har tillåtelse att satsa eller delta i aktiviteter, spel, programvara eller Speltjänster (även kollektivt häri kallat ”Tjänster”) på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] och [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], eller invånarna från USA eller Turkiet där tjänstera är stängt förbjudna.Om det kommer till[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]suppmärksamhet genom säkra källor att registrerade användare är en person under 18 år eller inte har rätt att använda Tjänstera, kommer [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], bland andra tillgängliga resurser, att avsluta den användarens konto. <br/>Detta avtal gäller till vilken använding som helst av Tjänsterna. I något fall av motstridelse mellan en bestämmelse av avtalet och någon bestämmelse på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]sPoker webbsida, företräder bestämmelsen av det här avtalet. Om inget häri motsäger det, med referens gjord i detta avtal till[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] ska anses ha gjorts till [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], och dess ansluta företag, efterträdare och övertagare. <br/>Dessa villkor, tillsammans med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Turnerings sektionen, Hur man spelar sektionen, alla spelregler, frånkopplingen och avslutningspolicy, och andra regler, policier och villkor på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] vilket specifikt relaterar to och styr vilka specifika händelser, spel, programvara eller turnering som helst utgör ett legalt bindande avtal (”Avtal”). Om detta avtal är översatt, ska den engelska texten ha företrädelse. Om något annat dokument ges i samband med detta avtal ska vara på engelska eller ska vara korrekt översatta på engelska och den engelska översättningen ska ha företrädelse i vilket fall som helst om några konflikter eller skillnader uppstår mellan dem. <br/><br/><strong>PROGRAMVARA</strong><br/><span style="font-weight: bold;">1.    LICENS FÖR PROGRAMVARA: </span><br/>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] bidrar en personlig, icke-exclusiv, icke överförbar licens att använda programvaran till dig, men behåller sig äganderätten till Programmvaran. Alla rättigheter som inte specifikt beviljas i detta avtal är reserverade av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] och, som tillämpade, [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s licensgivare. Mjukvaran är licenserad för ditt personliga bruk. Din licens ger ingen titel eller ägande i programvaran och ska inte tolkas som ett köp av några rättigheter i programvaran. <br/><br/><span style="font-weight: bold;">2.    ÄGANDE AV PROGRAMVARAN: </span><br/>Alla rättigheter, titlar och intressen och immateriella rättigheter till programmvaran ägs av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] eller dess licensgivare, och kan vara skyddade av tillämpade upphovsrätter eller andra immateriela rättigheter och spelregler och föredrag. Alla rättigheter som uttryckligen inte beviljats enligt detta avtal är reserverade av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].<br/><br/><span style="font-weight: bold;">3.    ANVÄNDNING AV PROGRAMVARAN: </span><br/> Du får endast använda programvaran i enighet med detta avtal. Du kan installera programvaran eller andra komponenter av tjänsterna på vilken annan personlig dator osm helst. Du kan göra säkerhetskopior av programvaran som ges då sådan användning och kopiering är för ditt personliga bruk i enighet med detta avtal, dessutom, sådana installationer och användningar görs endast via en dator där Du är den primära användaren. Du kan endast använda ett exemplar av programvaran på en dator åt gången. Du har inte tillåtelse att spela vid samma omgång eller i samma turnering med flera konton från samma hårdvara och genom att göra det bryter Du direkt mot detta avtal. <br/><br/><span style="font-weight: bold;">4.    BEGRÄNSNINGAR AV PROGRAMVARAN:</span><br/>Programvaran innehåller upphovsrättsskyddat material, affärshemligheter och annat egenutvecklat material. Du förstår att programvaran kodningsformat förblir en konfidentiell affärshemlighet av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Du får inte dekonstruera, dekompliera, modifiera, offentligt visa, förbereda härledda verk baserade på, ta isär eller på annat sätt reproducera eller ge andra möjlighet att använda programvaran. Du får inte sälja, tilldela, vidarelicensiera, hyra, låna ut eller direkt eller indirekt överföra programvaran till en tredje part. Varje handling i strid med detta avtal är oacceptabla.<br/><br/><span style="font-weight: bold;">5.    ÄNDRINGAR I FUNKTIONERNA AV PROGRAMVARAN: </span><br/> Genom att acceptera villkoren av detta avtal, går Du med på att[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] har tillåtelse att begränsa, neka, uppdatera eller avsluta några eller alla funktioner av denna programvara när som helst, utan några förvarningar. Du samtycker att bära riskerna av och hålla [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]menlös för några som helst ändringar och alla effekter av vad en ändring i fuktionerna kan påverka Din förmåga att använda programvaran.[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]kan kräva, som ett tillstånd, i din fortsätta tillgänglighet till[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]stjänster, accepterar Du att programvaran förbättras, justeras, anpassas, konverteringas till mer uppdaterade versioner av programvara eller att andra ändingar i programvara sker. <br/><br/><span style="font-weight: bold;">VILLKOR FÖR TJÄNSTERNA</span><br/><span style="font-weight: bold;">6.    ACCEPTERANDE AV VILLKOREN:</span><br/>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]tillåter Din användning av eller spelandet med dess tjänster, under förutsättning att Du följer villkoren av detta avtal. Vänligen läs dem noga. Genom att registrera och öppna ett konto som en kontemplation av sektion 7 nedan, försäkar Du att Du samtycker att hållas under villkoren av detta avtal. Om du inte vill vara bunden till dessa villkor, ska du inte registera dig och öppna ett konto, och Du kommer då inte få tillgång till eller använda tjänsterna. Villkoren för detta avtal kan ändras eller uppdateras när som helst av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)],utan att meddela Dig. Din fortsatta tillgång till, och användning av, tjänsterna kommer betyda att du samtycker att vara bunden till den mest uppdaterade versionen av detta avtal. Du kan se den mest uppdaterade verionen av detta avtal när som helst. <br/><br/><span style="font-weight: bold;">7.    REGISTRERING:</span><br/>För att använda [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]stjänster, måste Du först öppna ett konto genom att fylla i en unik och giltig e-mailadress och tillhörande lösenord. För att sätta in pengar på ditt konto måste du fylla i för- och efternamn, adress och telefonnummer. Du samtycker att förse endast sann och aktuell information och Du samtycker att uppdatera denna information när så är nödvändigt för att låta informationen förbli sann och uppdaterad. Du samtycker också till att låta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]sprogramvara ta ett digitalt fingeravtryck av din dator av säkerhetsskäl. Fingeravtrycket innefattar en uppsättning siffror, inklusive IP-konfiguration vilket sparas tillsammans med din information på kontot.När man öppnar ett konto med använding av riktiga pengar på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)],kommer Du kunna ha tillgång till följande: spela pengaspel, spela pengaspel turneringar. Med ett riktigt pengakonto, har Du tillgång till riktiga pengaspel och riktiga pengaturneringar. Det är strikt förbjudet att ha mer än ett aktivt konto på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] när som helst. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att stänga av, modifiera, ta bort och/eller lägga till några Spel med direkt verkan och utan att meddela Dig och[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]kommer inte vara ansvarig för sådana handlingar<br/><br/><span style="font-weight: bold;">8.    PERSONLIG ANVÄNDING AV SPELTJÄNSTERNA:</span><br/> Du samtycker att du håller din kontoinformation hemlig och konfidentiell och inte låta någon annan använda eller tillgå informationen. Allt deltagande i spel är Ditt val, och din risk. Genom att spela på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)],samtycker Du att Du inte kommer hitta Tjänster eller andra aspekter av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] som kan vara stötande, anstötande, orättvisa eller opassande. Du är endast tillåten att satsa för Din egen personliga underhållning. Andra kommersiella bruk av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] är förbjudet. Du samtycker att du är ansvarig för att kontrollera och följa lagarna som styr spel på den plats där programvaran används. <br/><br/><span style="font-weight: bold;">9.    ROBOTAR, ARTIFICIELLA INTELIGENSSYTEM OCH ANDRA SYSTEM:</span><br/>Det är högst förbjudet att använda några som helst automatiserade programvaror eller datorsystem för att spela på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)],inklusive agerandet att sända information från din dator till en annan dator där sådan programvara eller system är aktiverat. Poker robotar eller andra programvaror designade för att spela automatiskt på pokersidor är inte tillåtet. När än Du spelar på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)],kan programvaran skanna din dator för någon som helst aktivitet av ett sådant programvara eller system. Det är också förbjudet att använda någon typ av programvara under spelet som är designat för att spåra och visa handlingar från de andra spelarna på sidan eller andra system eller tjänster som överför medel till eller från en annan spelares[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto till deras konto på någon annan sida eller medvetet ”dumpa” av markörer mellan olika konton på CAKE poker nätverk. Använding av sådana metoder kommer resultera i att Ditt konto stängs av och dina vinster och pengar kommer konfiskeras. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att publicera information av något dokumenterat missbruk, inklusive Din personliga information.br/><br/><span style="font-weight: bold;">10.    INGA ANSTÄLLDA FRÅN FÖRETAGET:</span><br/>Om Du är en tjänsteman, direktör, anställd, konsult eller agent i Bolaget eller något av dess koncernbolag eller leverantörer eller försäljare, du är inte tillåtet att registrera sig med[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]eller delta varken direkt eller indirekt i några utav [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]sspeltjänster (som ”obehörig person”), om du gör så basserad på det skrivna tillåtandet av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]och sådant deltagande är en del av din anställning och/eller görs som marknadsföring för[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Släktingar med obehöriga personer har inte heller tillåtelse att registrera sig på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]eller delta varken direkt eller indirekt i några utav tjänsterna. I detta sammanhang syftar termen ”släkting” på (men inte endast begränsat till) make, sambo, förälder, barn eller syskon.<br/><br/><span style="font-weight: bold;">11.    SPELPENGAR:</span><br/>Spelpengar är inte riktiga (äkta) pengar och hålls separat från riktiga pengar. Spelpengar utgör inte eller representerar inte något värde alls. Spelpengar kan endast användas för att spela på bord där de använder spelpengar och kan inte samlas, betalas ut eller in på något annat sätt bli eller överföras mellan[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]och Dig eller någon annan person eller juridisk verksamhet.<br/><br/><span style="font-weight: bold;">12.    RIKTIGA PENGAR:</span><br/>För att spela med riktiga pengar, måste Du sätta in riktiga pengar på Ditt konto med någon utav metoderna som finns tillgängliga för dig från[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Minimala så väl som maximala gränser finns på överföringar av riktiga pengar. Alla äkta pengar kommer att betalas, spåras och behållas i US Dollar, och kommer inte ha någon ränta. Alla uttaxerade avgifter som betalas av processorer är Ditt ansvar. Genom att använda ditt kreditkort för att betala Ditt[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto kan behandlas som ett Cash Advance av banken som tar hand om ditt kreditkort. All ränta och/eller avgifter som associeras med ett Cash Advance är ditt ansvar. Vänligen se till att dina betalningar sker relativt snabbt. Om du betalar på mer än ett bord och [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] får för många klagomål gällande hastigheten på dina betalningar, kan[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]begränsa antalet bord du kan spela på samtidigt. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] är inte ansvarig för förluster som uppkommit på grund av oavsiktliga vad som sats av dig under ett spel eller när du spelar på flera bord och på grund av bord som byter plats på skärmen. Vänligen se till att du spelar på din skicklighetsnivå när du spelar på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].<br/><br/><span style="font-weight: bold;">13.    UTBETALNINGAR:</span><br/> I kassasektionen i programvaran kan du övervaka ditt saldo på kontot vilket är mängden riktiga pengar som du har tillgängliga, plus eller minus ackumulerade vinster eller förluster från att ha spelat några spel på Tjänsten, minus mängden som tidigare tagits ut av dig eller mängden pengar som förverkats eller återkrävts av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Alla pengar som tagits ut är en del mot transaktionsgränen och bearbetningsavgifter från [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Gränser och avgifter kan komma att ändras med tiden på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s egna initiativ eller av Dig ifall du anger specifika gränser. Utbetalningar utförs endast via metoderna som finns tillgängliga av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]i kassasektionen av programvaran och är, som standard, tillbakavisad med samma metod som föregående insättningar<br/><br/><br/><span style="font-weight: bold;">14.    SÄKERHETSKONTROLLER OCH FULLMAKTER:</span><br/>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att kontrollera Din identitet och trovärdigheten av informationen du har lämnat genom att göra olika säkerhet och ID-kontroller. Om Du misslyckas eller vägrar på företagets begäran och signerar en säkerhetsbegäran från[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], förbehåller[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sig rätten att ogiltigförklara ditt konto.<br/><br/><strong>15.</strong>    Om ingen överföring har registrerats på en spelares konto på 30 dagar, ska saldot på det kontot överföras till spelaren, eller om spelaren inte kan hittas, ska saldot överföras till LGA<br/><span style="font-weight: bold;"><br/>16.    [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] HÄNVISA-EN-VÄN PROGRAMMET:</span><br/>Genom att acceptera detta avtal, samtycker du att tillåta att[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] belönar Dig med bonusar med riktiga pengar för att du har hjälpt andra spelare att öppna ett riktigt pengakonto. Detta stöd materialiseras i allmänhet när du distribuerar din e-postadress till andra spelare och värvar dem genom att referera din e-postadress när de skapar ett konto.[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kan, ibland, erbjuda andra kampanjer eller initiativ designade för att assistera Dig med belöningar när du introducerar riktiga pengaspelare till [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] är inte ansvarig för misslyckandet av att en hänvisad spelare korrekt skickat hans/hennes e-mailadress.[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att ändra regler, nivåer och gränser på Hänvisa en vän programmet och dess riktning. <br/><br/><strong>17.</strong>    <br/>1.    Betalningar: Ditt konto kommer att få en bonus från Hänvisa en vän[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] programmet inom sju dagar från slutet på varje kalendermånad. <br/>2.    Att låsa upp nivåer och associerade bonusar: Regler styr hur man låser upp nivåer och de associerade bonusarna återfinns inuti [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s programvara. ( Klicka på Belöningar ->Hänvisa en Vän länken). Bonusar baseras på poäng från Frekventa spelare som genereras av spelarna Du har hänvisat. Om du misslyckas med att nå kraven för att få Frekventa Spelarpoäng på någon nivå, oavsett anledningen, kommer det resultera i att nivåerna förblir låsta eller outtagna.<br/>3.     Felaktig reklammetoder: Felaktig reklammetoder:[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]kommer belöna Dig om du berättar för andra om våra Speltjänster. Vi bevakar dock metoderna som används för att marknadsföra[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]och om det visar sig att du:<br/>4.    <br/>a.    Gör massutskick till oönskade e-postadresser<br/>b.     Medvetet och flagrant ignorera regler från någon 3:e parts webbplats genom att lägga inbjudningar att registrera sig, och/eller<br/>c.    Använder marknadsföringsmeddelande med grovt missledande påstående av PR belöningar<br/>Kan Du bli som deltagare få Ditt deltagande i [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]Hänvisa en vän programmet avbrytet eller avslutat. <br/><br/><br/><strong>18.</strong><br/>4.    Avslutandet av Hänvisa en vän deltagandet: Om utförandet av någon av de felaktiga reklammetoderna som beskrivs ovan utförs kan det resultera i din Uppsägning av deltagandet i Hänvisa en vän[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]programmet. Detta inkluderar en förlust av din nuvarande saldo från Hänvisa en vän programmet, förlust av framtida intäkter från Hänvisa en vän och borttagandet av förmågan för dig att hävda någon ytterligare hänvisade vänner.<br/><br/><span style="font-weight: bold;">19.    GULDKORT:</span><br/>Genom att acceptera detta avtal samtycker du att tillåta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] att belöna dig med Guldkort på ditt ringspel med riktiga pengar.I händelsen av att ett pris meddelas för ett Guldkort som du har för tillfället har du ansvaret att lösa Guldkortet före det offentliggjorda utgångsdatumet. Inget Guldkort kommer att tillåtas att lösas in mot ett pris när priset har gått ut. Ditt Guldkort kommer inte gå ut och kommer stanna på ditt konto, så länge kontot inte överges (se avsnitt 15).<br/><br/><span style="font-weight: bold;">20.    GULDMARKÖRER:</span><br/>Genom att acceptera detta avtal tillåter du [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] att belöna dig med Guldmarkörer baserat på reglerna som bestämts på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s webbsida). Din(a) Guldmarkör(er) kommer inte gå ut och kommer att stanna på Ditt konto, så länge kontot inte överges (se avsnitt 13).<br/><br/><span style="font-weight: bold;">21.   DRIFT AV DITT KONTO:</span><br/>Under villkoren för Ditt konto kan det uppkomma omständigheter som kräver ändrigar på Ditt konto. <br/><br/><strong>22.<br/></strong>1.    Succession: I händelse av Din död eller permanent inkapacitet, kräver[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]en kopia på dödscertifikatet eller en registrerad läkares medicinska utlåtande och alla andra handlingar som rör förvaltning eller förmyndarskap av din egendom som bevis på din efterträdare har eller vårdnadshavarens (gemensamt kallade "Förmånstagare") rätt. I denna händelse, kan dina inkomsträttigheter och/eller värdet av Ditt konto ges till Dina Förmånstagare. Dina förmånstagare måste skicka en skriven applikation styrkt av den nödvändiga dokumentationen som inkluderar dödscertifikatet eller en registrerad läkares medicinska utlåtande, för behandling av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].Godkännandet av denna applikation ska inte vara på orimliga grunder. Överföringar kommer endast godkännas om mottagarna är överens om att ta ansvar för Ditt konto dess skyldigheter som anges i dessa Villkor. Om mottagaren inte är tillåten att inneha ett konto, kommer bidragsmottagaren ha rätt att föra intresset av ditt konto till en tredje part som har rätt att inneha ett[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto. <br/>2.    Självutslutning: [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] förbehåller sig rätten att bevaka aktiviteten på ditt konto och meddela Dig om[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] tror att Du kan ha ett spelmissbruk. Hur som helst gör[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]inga garantier om dess förmåga att identifiera och hjälpa dig med spelmissbruk. Du kan begära att uteslutas från att komma in eller använda[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]stjänster av olika anledningar och du kan göra detta när som helst genom att skicka en begäran till <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br/>3.     Suspensioner och uppsägning av kontot:[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att avsluta Ditt konto när som helst om du bryter mot något av villkoren för Tjänster; eller ger falsk eller missledande information till[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)];eller tar del av bedrägligt, olämpligt eller stötande beteende mot[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] eller några andra av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s användare; eller är delaktiga i en aktivitet vilket kan anses strida mot vedertagna normer för god sed, i strid med tillämplig lagstiftning i Din juristdiktion och/eller strider mot intressena av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]eller som skadar[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s rykte. Sådana avslut ska göras av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]enligt eget gottfinnande men, handlingarna som kan uppkallas av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]i händelse av att du engagerar dig i sådant beteende kan inkludera, men är inte begränsade till varningar, tillfällig avstäningar av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s tjänster och, tillfällig avstäning av ditt[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto.<br/><br/>Avslutandet av ditt[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto kommer endast övervägas vid de allvarligaste överträdelserna eller som ett resultat av flera överträdelser och om möjligt endast efter upprepad kommunikation med dig. I händelse av uppsägning av ditt[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]konto ska[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]ha rätt att vidta sådana åtgärder som den anser lämpliga, inklusive att omedelbart blockera tillgången till[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s Speltjänster, beslagta alla pengar som finns på ditt konto med riktiga pengar, avslöjar sådan information (inklusive din identitet) till banker, kreditkortsföretag och/eller någon person eller enhet som har laglig rätt till sådan information, och/eller vidta rättsliga åtgärder mot dig. I händelse av uppsägning av ditt konto samtycker du:<br/>a.      till att Dina rättigheter att göra representationer gällande[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]som på något sätt omedelbart återkallas;<br/>b.       Dina rättigheter att använda[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s Tjänster, Ditt användarkonto och lösenord kommer omedelbart återkallas; <br/>c.       Du måste förstöra/ta bort alla Dina kopior av programvaran.<br/>d.       Dina rättigheter till eventuella befintliga eller framtida rättigheter Du annars kan ha haft eller har haft till följd av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]eller Din använding av[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)s tjänster, från och med dagen för uppsägning återkallas, och<br/>e.      Alla andra rättigheter under dessa Villkor och Tjänster är avslutade. <br/>4.    Restriktioner av chattande<br/>-    Du borde inte skriva om en hand medan den utvecklas.<br/>-    Du borde inte använda chatten för att erbjuda råd till andra spelare under en omgång, eller uppmana en spelare att göra en viss åtgärd.<br/>-    Du borde inte chatta om några som helst vikta kort du har haft på handen eller andra nuvarande kort du har på handen.<br/>-    Du borde endast chatta på engelska och bordets specifika språk som designats av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] för just det ändamålet.<br/>-     Du ska inte använda fula eller kränkande ord eller ett hotfullt språk.<br/> Ovanstående åtgärder motarbetas eftersom de visar dålig poker etikett och kan resultera i en suspension avchatten eller i svåra och kontinuerligt brytande fall ett komplett chattförbud eller stängning av konto.    <br/>5.     Andra brott mot någon del av dessa villkor för tjänster kan också resultera i förlust av någon eller alla befintliga krediter, arrende, priser eller vinster från spelverksamhet och alla andra rättigheter Du annars har eller har haft till följd av ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto eller Din använding av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s tjänster.[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] förbehåller sig också rätten att kräva ersättning för förluster till följd av bristande efterlevnad av de skyldigheter som följer av dessa användarvillkor. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] förbehåller sig rätten att stänga och avsluta Ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto för vilka välgrundade anledningar som helst när som helst utan att meddela dig.<br/><br/><span style="font-weight: bold;">23.     UTLÄMNANDE TILL TREDJE PART:</span><br/> Du samtycker till att hålla ditt konto och relaterad information hemlig och konfidentiell och att inte låta någon annan använda den. Om du avsiktligt eller oavsiktligt, direkt eller indirekt, avslöjar e-post och/eller lösenord till någon annan, och det resulterar i att en tredje part deltar i [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]s tjänster med Ditt e-mail och lösenord, kommer deltagandet vara ogiltigt, och Du kommer inte att återbetalas eventuella förluster på[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], oavsett huruvida tredje part har ditt samtycke eller inte. Bolaget skall inte krävas för att upprätthålla e-post eller lösenord om du tappar bort, glömmer eller blir av med dendata eller annars inte kan komma in på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] på grund av något annat än bolagets fel.<br/><br/><span style="font-weight: bold;">24.    SKADEERSÄTTNING:</span><br/> Du samtycker till att gottgöra, försvara och hålla[Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)], och dess moderbolag, dotterbolag, närstående bolag, tjänstemän, direktörer, aktieägare, anställda, agenter, licensgivare och samarbetspartners från alla anspråk , förluster, skulder, krav, skador, kostnader eller utgifter (inklusive rimliga advokatkostnader), som uppstår från eller hävdas av någon tredje part som på något sätt (a) Din användning av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]sTjänster, eller någon annan produkt, tjänst eller kampanj du erbjudits av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]; (b) anspråk på intrång i tredje parts immateriella rättigheter, (c) uppladdning, publicering, e-post, reproducera, överföra eller på annat sätt distribuera något innehåll eller annat material som du, eller (d) brott mot någon av dessa användarvillkor av dig eller alla användare av ditt konto med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] förbehåller sig rätten att ta det exklusiva försvaret och kontroll