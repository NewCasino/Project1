﻿Belopp som överförs till kort {0}
