﻿Januari