Välj konto för kreditering