Måndag