﻿Validation kod måste vara 6 tecken