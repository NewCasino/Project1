﻿An error has occurred during transaction processing.