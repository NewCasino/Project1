Välj en bonus