Ny e-mailadress