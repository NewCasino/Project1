﻿Ewire