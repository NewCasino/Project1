﻿Ditt namn här
