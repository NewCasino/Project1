Ange namnet på ditt konto