﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Ditt uttag-Ukash voucher
