Vänligen notera att det är olika begränsingar för maxbelopp gällande Ukash kort när det är utfärdat i en annan valuta. <table> <tr><td>Euro</td><td> : </td><td>EUR 250</td></tr> <tr><td>Australian Dollar</td><td> : </td><td>AUD 300</td></tr> <tr><td>Canadian Dollar</td><td> : </td><td>CAD 300</td></tr> <tr><td>Swiss Franks</td><td> : </td><td>CHF 300</td></tr> <tr><td>Czech Koruna</td><td> : </td><td>CZK 6000</td></tr> <tr><td>Danish Krone</td><td> : </td><td>DKK 1500</td></tr> <tr><td>Hungarian Forint</td><td> : </td><td>HUF 75000</td></tr> <tr><td>Latvian Lats</td><td> : </td><td>LVL 175</td></tr> <tr><td>Mexican Peso</td><td> : </td><td>MXN 4000</td></tr> <tr><td>Norwegian Krone</td><td> : </td><td>NOK 1500</td></tr> <tr><td>New Zealand Dollar</td><td> : </td><td>NZD 350</td></tr> <tr><td>Polish Zloty</td><td> : </td><td>PLN 1000</td></tr> <tr><td>Russian Ruble</td><td> : </td><td>RUB 9000</td></tr> <tr><td>Swedish Krone</td><td> : </td><td>SEK 2000</td></tr> <tr><td>US Dollar</td><td> : </td><td>USD 300</td></tr> <tr><td>South African Rand</td><td> : </td><td>ZAR 3000</td></tr> <tr><td>Sterling</td><td> : </td><td>GBP 200</td></tr> </table>