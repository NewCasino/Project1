﻿/game/gamerules.jsp?game=simsalabim&lang=sv