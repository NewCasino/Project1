<ol> <li><strong>INTRODUCTION:</strong><p>1.1.    By using and/or visiting any section of the website [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]   (the "Website"); or by opening an account on the Website you agree to be bound by:<br/>1.1.1.    the General Terms and Conditions, on this page; <br/>1.1.2.    the Privacy Policy,<br/>1.1.3.    any game rules,<br/>1.1.4.    any terms and conditions of  promotions, bonuses and special offers which may be found on the Website from time to time.<br/>1.2.    All of the terms and conditions listed above shall together be referred to as "the Terms".<br/>1.3.    Please read the Terms carefully before accepting them. If you do not agree to accept and be bound by the Terms please do not open an account or continue to use the Website. Your continued use of the Website constitutes acceptance of the Terms.<br/>1.4.    The Terms will come into effect on the 9th of June 2010.</p></li><li><strong>PARTIES</strong><p>2.1.    The Sportsbook Services and Content at the Website is provided by EveryMatrix Ltd, reg. no. C44411, 712, 14/19 Street, Valletta, VLT 1432 Malta. EveryMatrix maintains and operates a fully managed Sportsbook, by virtue of Letter of Intent Number LGA/CL2/497/2008 as issued by the Maltese Lotteries and Gaming Authority under the laws of Malta.<br/>2.2.    References in the Terms of Use to "us", "our," "we" or the “Company” are references to the party with whom you are contracting with, as specified above.</p></li><li><strong>CHANGES TO THE TERMS OF USE</strong><p>3.1.    We may need to change the Terms for a number of reasons, including for commercial reasons, to comply with new laws or regulations or for customer service reasons. The most up-to-date Terms of Use can be accessed here, and the date on which they came into force is noted.<br/>3.2.    Where we make changes to the Terms of Use which we wish to notify you of, we will do so by email or by placing a notice on the Website.</p></li><li><strong>OPENING YOUR ACCOUNT</strong><p>4.1.    In order to place a bet via the Website, you will need to open an account on the website ("Your Account").<br/>4.2.    For various legal or commercial reasons, we do not permit accounts to be opened by, or used from, customers based or domiciled in certain jurisdictions, including the United States of America. If you are in such a jurisdiction than you should not open an account or use the Website.<br/>4.3.    In order to open Your Account for use of the Website, You can contact Customer Services, or by clicking here and following the on-screen instructions.<br/>4.4.    When you open Your Account You will be asked to provide us with personal information, including your name, date of birth, and appropriate contact details, including an address, telephone number and e-mail address ("Your Contact Details"). <br/>4.5.    You hereby acknowledge and accept that, by using the services at the Website, you may both win and lose money.<br/>4.6.    Your Account must be registered in your own, correct, name. You may only open one account for the sportsbook. Any other accounts which you open with us in relation to the Service and the Website shall be "Duplicate Accounts". Any Duplicate Accounts may be closed by us immediately and:<br/>4.6.1.    all transactions made from the Duplicate Account will be made void;<br/>4.6.2.    all stakes or deposits made using that Duplicate Account will be returned to You; and<br/>4.6.3.    any returns, winnings or bonuses which you have gained or accrued during such time as the Duplicate Account was active will be forfeited by you and may be reclaimed by us, and you will return to us on demand any such funds which have been withdrawn from the Duplicate Account<br/>4.7.    If you wish to open another account, you may do so by contacting the Manager at <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>. If a new account is opened, the old account will be closed.<br/>4.8.    You must maintain your account and keep your details up-to-date.</p></li><li><strong>VERIFICATION OF YOUR IDENTITY; MONEY LAUNDERING REQUIREMENTS</strong><p>5.1.    You warrant that:<br/>5.1.1.    You are not younger than:<br/>5.1.1.1.    of 18 (eighteen) years; or<br/>5.1.1.2.    any legal age at which gambling or gaming activities under the law or jurisdiction that applies to you require ("the Legal Age"); and<br/>5.1.2.     the details supplied when opening Your Account are correct; and<br/>5.1.3.    You are the rightful owner of the money in your Account.<br/>5.2.    By agreeing to the Terms you authorise us to undertake verification checks as we may require ourselves or may be required by third parties (including, regulatory bodies) to confirm your identity and contact details (the "Checks"). <br/>5.3.    While we are undertaking any Checks, we may restrict you from withdrawing funds from Your Account. <br/>5.4.    In certain circumstances we may have to contact you and ask you to provide further information to us directly in order to complete the Checks. If you do not or cannot provide us with such information then we may suspend Your Account until you have provided us with such information or permanently close Your Account. Additionally, you will have to provide identification whenever you make a withdrawal of funds amounting to Two Thousand Three Hundred Euros (EUR 2,300) or more.<br/>5.5.    If we are unable to confirm that you are the Legal Age then we may suspend Your Account. If you are proven to have been under that age at the time you made any gambling or gaming transactions, then:<br/>5.5.1.    Your Account will be closed;<br/>5.5.2.    all transactions made while you were underage will be void, and all related funds deposited by you will be returned;<br/>5.5.3.    any stakes for bets made while you were underage will be returned to you; and<br/>5.5.4.    any winnings which you have accrued during such time will be forfeited by you and you will return to us any such funds which have been withdrawn from your Account.</p></li><li><strong>USERNAME, PASSWORD, AND CUSTOMER INFORMATION</strong><p>6.1.    After opening Your Account, you must not disclose (whether deliberately or accidentally) your username and password to anyone else. If you have lost or forgotten Your Account details you may retrieve your password by clicking on the “Forget your Password” link below the login portal.</p></li><li><strong>DEPOSITS AND WITHDRAWALS FROM YOUR ACCOUNT</strong><p>7.1.    If you wish to participate in betting or gaming using the Website, You must deposit money into Your Account which you can then use to place bets or play games. <br/>7.2.    Deposits to and withdrawals from an Account may be made through various payment providers that may change from time to time. Procedures, terms, and conditions vary between payment providers. We do not accept cash funds sent to us. <br/>7.3.    By depositing money you agree not to make any charge-backs, reversals or otherwise cancel any deposits into Your Account, and agree to refund and compensate us for unpaid deposits.<br/>7.4.    Your Account is not a bank account and is therefore not insured, guaranteed, sponsored or otherwise protected by any banking insurance system. Additionally any money deposited with us in your Account will not earn any interest. <br/>7.5.    We may at any time set off any positive balance on Your Account against any amount you owe to us when we re-settle any bets or wagers pursuant to Duplicate Accounts, Collusion, Cheating, Fraud and Criminal Activity or Errors.<br/>7.6.    You are responsible for reporting your winnings and losses to your local tax or other authorities.<br/>7.7.    You may request withdrawal of funds from Your Account at any time provided that:<br/>7.7.1.    all payments made into Your Account have been confirmed as cleared and none have been charged-back, reversed or otherwise cancelled;<br/>7.7.2.    any Checks referred to in paragraph 5 above have been completed. <br/>7.8.    Once we have approved your withdrawal you must give us sufficient information as to how the funds should be transferred to you. We will attempt to accommodate your request regarding the payment method and currency of your withdrawal. This, however, cannot be guaranteed. <br/>7.9.    We reserve the right to charge a fee amounting to our own costs (including the cost of the deposits) for withdrawals of funds that have not been put into play.<br/>7.10.1. Players who register with [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] must deposit from an account that is registered in their own name.<br/>7.10.2. We do not accept 3rd party deposits, ie. a friend, relative, partner, husband or wife.<br/>7.10.3. If we discover during our routine security checks that this has occurred, all casino winnings will be forfeited and sent back to the casino and the original deposit to the rightful owner of the account/Credit Card.<br/>7.10.4. If bank transfer is required to return the money to the rightful owner, all bank charges will be borne by the receiver.<br/>7.10.5. In case of mastercard deposits where refunds are not possible, The card owner must sign ‘credit card verification form’ and send in identification documents for us to do the verification.</p></li><li><strong>PLACING A BET OR GAMING</strong><p>8.1.    All transactions will be concluded in the language from which you placed your transaction.<br/>8.2.     It is your responsibility to ensure that the details of any transaction are correct. <br/>8.3.    You can access your transaction history on the Website.<br/>8.4.    We reserve the right to refuse the whole or part of any transaction requested by you at any time in our sole discretion. No transaction is accepted by us until we have confirmed to you that it has been accepted. If you do not receive a confirmation that your transaction has been accepted, you should contact Customer Services.<br/>8.5.    Once your bet is confirmed, you cannot cancel the transaction without our written consent.</p></li><li><strong>COLLUSION, CHEATING, FRAUD AND CRIMINAL ACTIVITY</strong><p>9.1.    The following activities as not allowed and constitute a material breach of the Terms: <ul> <li>colluding with other third parties; </li> <li>using unfair advantage or influence (commonly known as cheating), including the exploitation of a fault, loophole or error in our software, the use of automated players (sometimes known as 'bots'); or the exploitation of an 'error';</li> <li>undertaking fraudulent activities to your advantage, including the use of a stolen, cloned or otherwise unauthorised credit or debit card, as a source of funds;</li> <li>taking part in any criminal activities including money laundering and any offence with criminal repercussions.</li> </ul>9.2.    We will take all reasonable steps to prevent such activities; detect them and the relevant players; and deal with the relevant players appropriately. We will not be liable for any loss or damage which you or any other player may incur as a result of collusive, fraudulent or otherwise illegal activity, or cheating, and any action we take in respect of the same will be at our sole discretion.<br/>9.3.    If you suspect a person is colluding, cheating or undertaking a fraudulent activity, you shall as soon as reasonably practicable report it to us by e-mailing us.<br/>9.4.    We reserve the right to inform relevant authorities, other online gaming or gambling operators, other online service providers and banks, credit card companies, electronic payment providers or other financial institutions of your identity and of any suspected unlawful, fraudulent or improper activity, and you agree to cooperate fully with us to investigate any such activity.</p></li><li><strong>OTHER PROHIBITED ACTIVITES</strong><p>10.1.    You should not use the Website for any purpose which is considered to be defamatory, abusive, obscene, racist, sexist, discriminatory, or offensive. You must not use any abusive or aggressive language or images; swear, threaten, harass or abuse any other person, including other users, or behave in such a manner towards any Company staff used to provide the Website or Customer Services.<br/>10.2.    You shall not corrupt the Website, flood the Website with information so as to cause the Website to not function, nor use any features which may affect the function of the Website in any way for example (but not limited to) releasing or propagating viruses, worms, logic bombs or similar. Any multiple submissions or "spam" are strictly prohibited. You must not interfere or tamper with, remove or otherwise alter in any way, any information in any form which is included on the Website.<br/>10.3.    You shall use the Website for personal entertainment only and shall not be allowed to reproduce the Website or any part of it in any form whatsoever without our express consent.<br/>10.4.    You must not attempt to gain unauthorised access to the Website, the servers on which the Website is stored or any server, computer or database connected to the Website. You must not attack the Website via a denial-of-service attack or similar. When breaching this provision we will report any such breach to the relevant law enforcement authorities and we will co-operate with those authorities by disclosing your identity to them. In the event of such a breach, your right to use the Website will cease immediately.<br/>10.5.    We will not be liable for any loss or damage caused by a distributed denial-of-service attack, viruses or other technologically harmful material that may infect Your computer equipment, computer programs, data or other proprietary material due to Your use of the Website or to Your downloading of any material posted on such Website, or on any website linked to the Website.<br/>10.6.    It is prohibited to sell or transfer accounts between players.</p></li><li><strong>CLOSURE AND TERMINATION BY US</strong><p>11.1.    It is company policy in the interests of security and in accordance with Maltese legislation, that if no transaction has been recorded on Your Account for thirty months (an “Inactive Account”), we shall remit the balance in that account to you. If you cannot be satisfactorily located any funds in that account will be handed over to the Lotteries & Gaming Authority of Malta. Thus the funds are available to the player wishing to withdraw them.<br/>11.2.    Your Inactive Account will be terminated with written notice (or attempted notice) using your contact details. In the event of any such termination by us, other than where such closure and termination is made pursuant to paragraph 11 (Collusion, Cheating, Fraud and Criminal Activity) or paragraph 20 (Breach of the Terms of Use) of these Terms, we will refund the balance of Your Account to you. If you cannot be located, the funds shall be remitted to the relevant gambling authority. </p></li><li><strong>ALTERATION OF THE WEBSITE</strong><p>12.1.    We may, in our absolute discretion, alter or amend any product offered via the Website at any time for the purpose of maintaining the Website.  </p></li><li><strong>IT FAILURE</strong><p>13.1.    Where unexpected system flaws, faults or errors occur in the software or hardware which we use to provide the Website we will take immediate steps to remedy the problem. <br/>13.2.    We do not accept any liability for IT failures which are caused by your equipment used to access the Website or faults which relate to your internet service provider.</p></li><li><strong>ERRORS OR OMISSIONS</strong><p>14.1.    A number of circumstances may arise where a bet is accepted, or a payment is made, by us in Error. <br/>14.2.    [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] reserves the right to cancel any bet made on obviously incorrect odds, switched odds (where odds were listed against the wrong teams) or a bet made after an event has started if that event is not available for live betting. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] reserves the right to refuse, restrict, cancel or limit any bet.<br/>14.3.    Neither we (including our employees or agents) nor our partners or suppliers shall be liable for any loss including loss of winnings that results from any Error by us or an error by you. You will forfeit any winnings/losses that result from any such Error.</p></li><li><strong>EXCLUSION OF OUR LIABILITY</strong><p>15.1.    Your access to and use of the products offered via the Website, is at your sole option, discretion and risk. <br/>15.2.    We will provide the Website with reasonable skill and care and substantially as described in the Terms. We do not make any other promises or warranties the Website, or the products offered via the Website, and hereby exclude (to the extent permitted by law) all implied warranties in respect of the same.<br/>15.3.    We shall not be liable to You in contract, tort (including negligence) or otherwise for any business losses, including but not limited to loss of data, profits, revenue, business, opportunity, goodwill, reputation or business interruption or for any losses which are not currently foreseeable by us arising out of the Terms of Use or Your use of the Website.</p></li><li><strong>BREACH OF THE TERMS OF USE</strong><p>16.1.     You shall compensate us in full for any claims, liabilities, costs, expenses (including legal fees) and any other charges that may arise as a result of your breach of the Terms.<br/>16.2.    Where you are in material breach of the Terms, we reserve the right, but shall not be required, to:<br/>16.2.1.    Provide you with notice (using Your Contact Details) that you are in breach requiring you to stop the relevant act or failure to act,<br/>16.2.2.    suspend your Account so that you are unable to place bets or play games on the Website, <br/>16.2.3.     close Your Account with or without prior notice from us.<br/>16.2.4.    recover from Your Account the amount of any pay-outs, bonuses or winnings which have been affected by any material breach.<br/>16.3.    We have the right to disable any user identification code or password if in our reasonable opinion you have failed to comply with any of the provisions of the Terms.</p></li><li><strong>INTELLECTUAL PROPERTY RIGHTS</strong><p>17.1.    All website design, text, graphics, music, sound, photographs, video, the selection and arrangement thereof, software compilations, underlying source code, software and all other material contained within the Website are subject to copyright and other proprietary rights which are either owned by us or used under licence from third party rights owners. To the extent that any material contained on the Website may be downloaded or printed then such material may be downloaded to a single personal computer only and hard copy portions may be printed solely for your own personal and non-commercial use.<br/>17.2.     Under no circumstances shall the use of the Website grant to any user any interest in any intellectual property rights (for example copyright, know-how or trade marks) owned by us or by any third party whatsoever.<br/>17.3.    No rights whatsoever are granted to use or reproduce any trade names, trade marks or logos which appear on the Website except as specifically permitted in accordance with the Terms of Use.</p></li><li><strong>YOUR PERSONAL INFORMATION</strong><p>18.1.    We are required by law to comply with data protection requirements in the way in which we use any personal information collected from you in your use of the Website. We therefore take very seriously our obligations in relation to the way in which we use your personal information.<br/>18.2.    By providing us with the information, you consent to our processing your personal Information for the purposes set out in the Term, for operating the Website or to comply with a legal or regulatory obligation.<br/>18.3.    As a policy the Company will not disclose any personal information to anyone other than those employees that need access to your data to provide you with a service.<br/>18.4.    We will retain copies of any communications that you send to us (including copies of any emails) in order to maintain accurate records of the information that we have received from you.</p></li><li><strong>USE OF COOKIES ON THE WEBSITE</strong><p>19.1.    The Website uses 'cookies' to assist the functionality of the Website. A cookie is a small file of text which is downloaded onto your computer when you access the Website and it allows us to recognise when you come back to the Website. Information on deleting or controlling cookies is available at www.aboutcookies.org. Please note that by deleting our cookies or disabling future cookies you may not be able to access certain areas or features of the Website.</p></li><li><strong>COMPLAINTS AND NOTICES</strong><p>20.1.    If You wish to make a complaint regarding the Website, a first step should be to, soon as reasonably possible, contact Customer Services.<br/>20.2.    In the event of any dispute, you agree that the records of the server shall act as the final authority in determining the outcome of any claim.<br/>20.3.    You agree that in the unlikely event of a disagreement between the result that appears on your screen and the game server, the result that appears on the game server will prevail, and you acknowledge and agree that our records will be the final authority in determining the terms and circumstances of your participation in the relevant online gaming activity and the results of this participation.<br/>20.4.    When we wish to contact you regarding such a dispute, we will do so by using any of Your Contact Details.</p></li><li><strong>INTERPRETATION</strong><p>21.1.    The original text of the Terms is in English and any interpretation of them will be based on the original English text. If the Terms of Use or any documents or notices related to them are translated into any other language, the original English version will prevail.</p></li><li><strong>TRANSFER OF RIGHTS AND OBLIGATIONS</strong><p>22.1.    We reserve the right to transfer, assign, sublicense or pledge the Terms, in whole or in part, to any person, provided that any such assignment will be on the same terms or terms that are no less advantageous to You. </p></li><li><strong>EVENTS OUTSIDE OUR CONTROL</strong><p>23.1.     We will not be liable or responsible for any failure to perform, or delay in performance of, any of our obligations under the Terms of Use that is caused by events outside our reasonable control, including, without limitation, acts of God, war, civil commotion, interruption in public communications networks or services, industrial dispute or DDOS-attacks and similar Internet attacks having an adverse effect ("Force Majeure"). Our performance is deemed to be suspended for the period that the Force Majeure Event continues, and we will have an extension of time for performance for the duration of that period. We will use our reasonable endeavours to bring the Force Majeure Event to a close or to find a solution by which our obligations may be performed despite the Force Majeure Event.</p></li><li><strong>WAIVER</strong><p>24.1.    If we fail to insist upon strict performance of any of your obligations or if we fail to exercise any of the rights or remedies to which we are entitled, this shall not constitute a waiver of such rights or remedies and shall not relieve you from compliance with such obligations.<br/>24.2.    A waiver by us of any default shall not constitute a waiver of any subsequent default. No waiver by us of any of the provisions of the Terms shall be effective unless it is expressly stated to be a waiver and is communicated to you in writing in accordance with above.</p></li><li><strong>SEVERABILITY</strong><p>25.1.    If any of the Terms are determined to be invalid, unlawful or unenforceable to any extent, such term, condition or provision will to that extent be severed from the remaining terms, conditions and provisions which will continue to be valid to the fullest extent permitted by law. In such cases, the part deemed invalid or unenforceable shall be amended in a manner consistent with the applicable law to reflect, as closely as possible, Our original intent.</p></li><li><strong>LAW AND JURISDICTION</strong><p>26.1.    The Terms of Use shall be governed by and interpreted in accordance with the laws of England and Wales save for any issues arising in respect to the Maltese licence which will be governed by Maltese Law in the Maltese Courts.<br/>26.2.    The Courts of England and Wales shall have non-exclusive jurisdiction over any disputes arising out of the Terms of Use themselves.</p></li><li><strong>RESPONSIBLE GAMING AND GAMBLING</strong><p>27.1.    For those customers who wish to restrict their gambling, we provide a voluntary self-exclusion policy, which enables you to close Your Account or restrict your ability to place bets. If you require any information relating to this facility please speak to Customer Services.<br/>27.2.    We will use our reasonable endeavours to ensure compliance with your self-exclusion. However you accept that we have no responsibility or liability whatsoever if you continue gambling and/or seek to use the Website and we fail to recognise or determine that.<br/>27.3.    We are committed to supporting Responsible Gambling initiatives and encourage you to find information about Responsible Gambling at the websites of the following organisations:<br/>Gambling Therapy - www.gamblingtherapy.org<br/>Gordon House Association - <a href="http://www.gordonhouse.org.uk">www.gordonhouse.org.uk</a></p></li><li><strong>LINKS</strong><p>28.1.    Where we provide hyperlinks to other websites, we do so for information purposes only. You use any such links at your own risk and we accept no responsibility for the content or use of such websites, or for the information contained on them.</p></li> </ol><p style="text-align:right"> <button type="button" onclick="window.print(); return false" class="button"> <span class="button_Right"> <span class="button_Left"> <span class="button_Center"> <span>Print</span> </span> </span> </span> </button></p>