Skicka allt