﻿Nedtrappning under 3 månader
