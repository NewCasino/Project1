﻿Ange ett lösenord här
