För att bjuda in dina vänner till MamaPortal, skicka nedanstående länk till dem via e-post, IM, skype, etc.: