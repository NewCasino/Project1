﻿Sätt en insättningsgräns
