Klicka  <a href="http://www.smscoins.net" target="_blank">here</a> för att köpa mynt. 