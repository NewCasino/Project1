﻿Registrera Dig
