﻿Neteller(Ryssland)
