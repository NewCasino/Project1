﻿Välj Konto
