februari