﻿{0}m sedan