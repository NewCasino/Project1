﻿Macedonia