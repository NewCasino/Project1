Inget förfallodatum