Min favoritställe?