﻿Europeisk Roulette
