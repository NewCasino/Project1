Om du inte mottar ett e-postmeddelande inom kort, kontrollera din skräppostkorg.