﻿Tecken