﻿Lösenord:
