Endast siffror och punkt är tillåtna. Använd punkt som decimaltecken och ange oformaterad siffra.