﻿Nej
