Generera en kod för att kunna göra uttag från Bank of Georgias bankomat.