﻿Smeknamn
