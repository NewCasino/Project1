﻿Begränsningstyp
