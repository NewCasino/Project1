Ange lösenord