﻿Moneybookers-konto(n)
