1 års självuteslutningsperiod