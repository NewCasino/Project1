Ange kortnummer.