﻿User is not assigned the role '{0}'