﻿MasterCard