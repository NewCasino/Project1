Om inte mailet kommer fram inom några minuter, vänligen kolla skräp/spam korgen