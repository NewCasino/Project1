﻿Vänligen skriv in BIC
