Banköverföring online