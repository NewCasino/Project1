﻿Alla