Spela 