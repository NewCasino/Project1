Du har inga pågående uttag just nu. 
<br /><br />
När du har ett pågående uttag i listan nedan, har du möjlighet att avbryta den transaktionen och omedelbart föra tillbaka pengarna till ditt konto.