Du måste aktivera ditt konto först innan du kan spela i riktiga pengar-läge!