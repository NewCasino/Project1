Ditt namn