Plånbok nummer