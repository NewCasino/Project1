﻿Min antal poäng att växla in
