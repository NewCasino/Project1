Tjeckien, Koruny