Detta alias är inte tillgängligt eller används redan av andra, var vänlig försök med ett annat alias.