﻿Få exklusiva erbjudanden via SMS.
