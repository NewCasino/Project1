Spela LIVE Roulette nu!