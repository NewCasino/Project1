﻿Laddar Saldon
