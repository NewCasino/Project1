﻿Virgin Islands (U.S.)