Välj giltighetstid fr.o.m.