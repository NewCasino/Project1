﻿Registrera ett kort
