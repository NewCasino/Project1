﻿Trappa ned till
