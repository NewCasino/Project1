﻿Beloppet överskrider din dagliga gräns
