﻿Adress
