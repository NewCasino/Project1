﻿Växla
