﻿Oktober