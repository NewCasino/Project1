E-mailadress domänen är inte tillåten