﻿/game/gamerules.jsp?game=deuceswild5&lang=sv