﻿Uppfriska Balansen
