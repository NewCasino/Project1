Senaste bankkonton