﻿/game/gamerules.jsp?game=krakow&lang=sv