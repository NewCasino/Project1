Ange ditt ID-nummer