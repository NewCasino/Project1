Lyckad