﻿Överföring till vän ej tillåten!
