﻿Belopp som satts in på ditt {0} konto