﻿You have requested an amount over EUR 2300, it is our legal requirement to verify you.Please send the following documents to support <br />
1. passport copy <br />
2, prove of address (utility bill or bank statement, less tha 3 month old) <br />
We will process the transaction after we have verified you