Användarnamnet måste bestå av minst 4 tecken