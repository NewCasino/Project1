Logga ut