﻿Uttag av pengar direkt till din bank via Intelligent Payments