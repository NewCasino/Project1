Ukash-värde