﻿Vänligen ange ditt UIPAS Konto ID.
