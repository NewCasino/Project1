﻿Max beloppet måste vara ett nummer.


