﻿vänligen ange en beskrivning
