Se föregående jackpot