﻿Tyvärr, din begäran om insättning {0} har nekats.<br />
Din bank kan ha restriktioner för hur ditt kort används online.<br /><br />
<strong>Våra föredragna betalningsalternativ: EntroPay!</strong><br />
Det är ett alternativt sätt att betala och som gör din insättning {1} 
lika enkel som 1-2-3!