Belopp som debiterats från ditt {0} konto