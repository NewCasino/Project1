Georgian Card- leverantörer för korthanterings tjänster