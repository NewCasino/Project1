﻿Du spelar med låtsaspengar.Logga in för att spela med riktiga pengar.
