﻿Upprepa ditt nya lösenord här

