Ange referensnumret.