Välj valuta