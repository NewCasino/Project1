﻿/game/gamerules.jsp?game=jokerwild25&lang=sv