Ditt förnamn måste innehålla minst 2 tecken