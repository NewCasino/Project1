Jag är {0} år eller äldre.