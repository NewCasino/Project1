Att sätta in på {0} konto