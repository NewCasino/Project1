﻿Uttag ej tillåtna!
