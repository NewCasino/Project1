Ogiltigt datum