﻿            <li class="GLItem BannerGLItem hidden">
                <a href="#" class="GameThumb BannerThumb" title="BannerThumb">
                    <span class="GameThumbContent">
                        <span class="GameBannerTitle">Turkish tables</span>
                        <span class="GameBannerSubTitle">online hours</span>
                        <span class="GameBannerDays">Monday,Wensday,Friday</span>
                        <span class="GameBannerHours">10:00am - 7:00pm</span>
                    </span>
                </a>
            </li>
