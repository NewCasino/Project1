Klassificering: