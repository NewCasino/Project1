﻿Din session har gått ut, vänligen logga in igen.
