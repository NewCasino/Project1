﻿Svenska kronor (SEK)