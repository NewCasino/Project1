Uttag till