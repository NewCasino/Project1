Tiden för den här sessionen har löpt ut, logga in igen.