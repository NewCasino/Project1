﻿<img src="//cdn.everymatrix.com/Shared/_files/Deposit/CardGuide_IssueNumber.png" />
<br />
<span>Om ditt kort saknar utgivningsnummer, lämna fältet tomt.  </span>