﻿Av säkerhetsskäl ber vi dig att ändra ditt lösenord så att lösenordet följer licensieringsreglerna.

