Min favorit seriefigur?