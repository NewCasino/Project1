Vänligen besvara säkerhetsfrågan