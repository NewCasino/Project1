﻿/game/gamerules.jsp?game=frog&lang=sv