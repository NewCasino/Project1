﻿<ol>
        
<li> <strong> Jag har laddat ner programmet - där är det </strong>?
<p> När [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] Pokers mjukvara har installerats på datorn, en [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] Poker-ikonen visas på skrivbordet. Helt enkelt dubbelklicka på den här ikonen för att starta pokerklienten och du ska tas omedelbart till vår Spellobby. </P>
</li>


<li> <strong> Min lösenordet inte accepteras? </strong>
<p> Ange ett felaktigt lösenord kan ofta resultera i en "inte kan validera lösenord" kod. Eftersom lösenord är skiftlägeskänsliga, kontrollera din Caps Lock är avstängd. Om dina problem kvarstår, välj "glömt lösenord"-knappen och ett nytt lösenord kommer att utfärdas till den e-postadress som anges på [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)]. Konto </p>
</li>


<li> <strong> Kan jag ändra mitt smeknamn? </strong>
<p> [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] Poker tillåter spelare möjligheten att ändra sitt spelar-ID (namn uppträder vid pokerborden) var 7 dagar. För att göra detta, besök "Mitt konto" när du är inloggad på den [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] Poker programvara </p>.
</li>


</ol>

<p style="text-align:right">
     <button type="button" onclick="window.print(); avkastning false" class="button">
         <span class="button_Right">
             <span class="button_Left">
                 <span class="button_Center">
                     <span> Print </span>
                 </span>
             </span>
         </span>
     </knappen>
</p>
