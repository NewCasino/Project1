Snabbregistrering