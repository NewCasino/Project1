Ditt förnamn måste bestå av minst 2 tecken