﻿/game/gamerules.jsp?game=kenobnjp&lang=sv