Förverkad