Australien Dollar