Din kompis användarnamn eller e-postadress är felaktig.