Tillåt mig inte att logga in någonsin igen