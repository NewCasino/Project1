﻿visa menyn
