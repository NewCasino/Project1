Vänligen fyll i bonusinehåll på/Metadata/Documents/NetEntTermsAndConditions.DefaultHtml