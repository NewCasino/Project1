Upprepa lösenordet