Online: