﻿/game/gamerules.jsp?game=hotcity&lang=sv