﻿Registrering öppen
