Visning