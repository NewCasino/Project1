Överföring