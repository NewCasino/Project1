Uttag av pengar direkt till ditt Voucher-konto