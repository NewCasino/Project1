Du måste logga in för att bjuda in en vän.