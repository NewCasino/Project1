Tyvärr, din aktivitet misslyckades, försök igen.