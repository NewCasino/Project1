﻿<img src="//cdn.everymatrix.com/_casino/1/1187C99038E5432A254DA3803941BF3A.jpg" />
