Insättning till