Gräns för negativt saldo