Kortets säkerhetskod (CVC)