﻿/game/gamerules.jsp?game=hilo&lang=sv