﻿[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Sport
