Konfiskera alla medel vid förverkande