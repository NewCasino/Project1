﻿Fröken