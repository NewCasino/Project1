﻿All American -sarja
