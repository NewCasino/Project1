﻿Franska Roulette Serier
