Ange mottagarens telefonnummer.