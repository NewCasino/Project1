﻿Banköverföring
