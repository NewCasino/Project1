﻿IGT
