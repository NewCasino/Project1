﻿EPS