Lokal bank