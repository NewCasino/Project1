En 7 dagars avstängning kan bara användas två(2) gånger