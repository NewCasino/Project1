Vänligen ange din email adress