Vänligen fyll kortets säkerhetskod.