﻿/game/gamerules.jsp?game=bloodsuckers&lang=sv