Populära spel