Problem med webbsidan