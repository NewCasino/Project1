﻿Inloggningen misslyckades. Ditt konto är på en nedtrappningsperiod som kommer utlöpa den {0}, försök logga in igen efter detta datum.
