﻿Alla Spel
