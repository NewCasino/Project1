﻿/game/gamerules.jsp?game=deuceswild25&lang=sv