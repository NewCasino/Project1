﻿Satsa på vår Odds
