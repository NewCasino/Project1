﻿<ol>
 <li> <strong>Hur öppnar jag ett [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto?</strong> 
 <p>**Du kan skapa ett konto [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] på något av följande sätt: 1)
 <a href="/regist>Klicka direkt här.</a>
 2) Eller så kan du gå till hemsidan och klicka på "Registrera" överst i vänstra hörnet eller på "Gå med nu" överst till höger. Oavsett vilket du väljer, kommer du att dirigeras till registreringssidan. Observera att ditt användarnamn och din kontovaluta inte kan ändras senare.
 <br />
Du kan även ange en kampanjkod. Innan du skickar dina uppgifter, se till att du försäkrar att du är över 18 år och godkänner våra "Villkor och bestämmelser". Du kan logga in på ditt konto direkt från valfri [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sida med hjälp av ditt användarnamn och lösenord.
 </p>
 </li>

 <li> <strong>Varför kan jag inte skapa ett konto?</strong>
 <p>
Kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kundtjänst på
 <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">
 [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]
 </a>
 så hjälper vi dig.
 </p>
 </li>

 <li>
 <strong>Varför måste jag skapa ett konto för att spela era spel?</strong>
 <p>
Vi vill att du öppnar ett konto [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] för att då godkänner och följer du våra regler och&nbsp; bestämmelser, som inkluderar en försäkran om att du är över 18 år.
 </p>
 </li>

 <li>
 <strong>Varför behövs mina personliga uppgifter? Är mina personliga uppgifter säkra hos er?</strong> 
 <p>
Vi behöver dina personliga uppgifter för att bekräfta din identitet, ålder, adressbevis och alla ekonomiska transaktioner.&nbsp; [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] använder de allra senaste datakrypteringsteknikerna för att skydda dina personliga uppgifter.
 </p>
 </li>

 <li>
 <strong>
 Måste jag göra en insättning för att kunna öppna ett konto hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]?
 </strong>
 <p>
 Nej, du kan spela i vårt Casino och spela Poker på skoj om du vill.
 </p>
 </li>

 <li>
 <strong>Kan jag ha mer än ett konto?</strong>
 <p>Nej, endast ett konto är tillåtet.</p>
 </li>

 <li>
 <strong>
 Finns det någon lägsta åldersgräns för att spela på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]?
 </strong>
 <p>
 Du måste vara minst 18 år för att spela på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sajten.
 </p>
 </li>

 <li>
 <strong>Accepterar ni spelare som är bosatta i mitt land?</strong>
 <p>
 Så länge du inte bryter mot några lagar i ditt land accepterar vi spelare från alla länder utom USA, Frankrike och Turkiet.
 </p>
 </li>

</ol>

<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Print</span>
 </span>
 </span>
 </span>
 </button>
</p>