Prova våra mini-spel!