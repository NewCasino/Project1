Login misslyckades.Kontrollera användarnamnet och lösenordet.