Uppdatera mobil