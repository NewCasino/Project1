﻿Spela i vårt Kasino
