Adressrad 1