﻿/game/gamerules.jsp?game=jacksorbetter5&lang=sv