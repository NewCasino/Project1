<p>Kära $USERNAME$, <br /><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Det här e-mailet bekräftar att du har ändrat din personliga tidsbegränsningar från $LIMITPERIOD$ minuter till $NEWLIMITPERIOD$ minuter. Den nya gränsen kommer att bli aktiverad på $LIMITEXPIRYDATE$. <br /><br /> Vänligen tveka inte att kontakta oss om du har några frågor på<ahref="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p><br /> Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>