﻿Ditt kumulativa uttag har överskridit 2300 EUR, enligt bestämmelser är vi tvungna att verifiera ditt konto innan vi kan bearbeta ditt uttag. Vänligen skicka ett E-post med följande dokument. <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>
<p>a) bevis på adress, till exempel faktura eller kontoutdrag </p>
<p>b) en kopia av ett nationellt ID eller pass</p>
<p>c) en kopia av kortet som användes vid insättning </p>



