Ogiltig kampanjkod.