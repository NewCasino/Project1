Skicka om verifieringskod