﻿Meddelandenummer till mottagare(Refcode)

