Meddelande till mottagare (Ref-kod)