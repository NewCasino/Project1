Ange ditt bankkontonummer