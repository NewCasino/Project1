﻿Kontaktuppgifter
