Spara