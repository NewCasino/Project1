﻿Vänligen skriv in din plånbok
