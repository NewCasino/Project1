﻿Daglig gräns
