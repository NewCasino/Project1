﻿Föregående sida
