﻿Starttid
