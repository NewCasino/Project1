Decimaler som inte är 0 accepteras inte av TLNakit