﻿Hjälp
