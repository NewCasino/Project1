Transaktionen är oavslutad, vänligen uppdatera denna sida efter avslutad transaktion.