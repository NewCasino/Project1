﻿AU$ (AUD)