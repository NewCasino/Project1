Var god och välj ett lösenord