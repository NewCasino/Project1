För att sättas in på {0} konto