﻿Vi ber om ursäkt men du är inte berättigad för överföring just nu. Vänligen <a href="/KontaktaOss">kontakta supporten</a> för mer information 
