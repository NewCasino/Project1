Ogiltig affiliate-markering i din url, vänligen kontrollera. 