Visa bord