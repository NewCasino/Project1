Gå med nu!