﻿/Casino/Info/fpp-räntesats
