﻿Välkommen till [Metadata:value(/Metadata/Settings.Operator_DisplayName)]
