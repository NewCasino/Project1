Uttag direkt till ditt ABAQOOS konto