Slutdatum måste infalla efter startdatum.