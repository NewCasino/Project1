Logga in först.