Föregående spel