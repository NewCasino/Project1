Bankkontots valuta