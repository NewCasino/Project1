Besök LIVE Casino lobbyn