Uttag av pengar direkt till ditt PaySafeCard-konto