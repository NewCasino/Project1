﻿<p class="ATHP">Tappa på <span class="ATHIcon">Lägg till hemskärm </span> ikonen nedan och välj "Lägga till hemskärm".</p>
