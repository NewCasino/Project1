﻿<p>Kära&#160; $USERNAME$,<br />
<br />
Tack för att du registrerat dig på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]
<br />
<br />
För din egen säkerhet vill vi påminna dig om att verifiera din e-postadress för att säkerställa att kontot förblir aktivt så att du kan fortsätta dra nytta av alla suveräna erbjudanden på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].<br />
<br />
Klicka på länken nedan, om den inte fungerar, försök kopiera och klistra in länken i din webbläsare.<br />
<br />
<a href="$ACTIVELINK$">$ACTIVELINK$</a></p>
<br />
Om du inte har registrerat dig hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]
, bortse från det här e-postmeddelandet eller meddela <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br />
<br />
Se till att slutföra din e-postverifiering direkt så att ditt konto inte blir begränsat för din säkerhets skull.
<p><br />
Vänliga hälsningar,<br />
[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]
 Kundtjänstteamet<br />