﻿Pöytäpelit

