﻿User is already assigned the role '{0}'