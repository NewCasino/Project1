﻿Voucher-nummer