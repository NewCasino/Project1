Se nästa jackpot