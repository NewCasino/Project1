Ange ett mobilnummer som innehåller mellan 7 -30 nummer