﻿Klicka för detaljer
