Visa {0}