﻿Vänligen välj kortet.
