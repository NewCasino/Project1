﻿Videokolikkopelit
