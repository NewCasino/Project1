Uttag av pengar direkt till ditt UseMyServices-konto