﻿<ol>

 <li> <strong>Hur gör jag en insättning på mitt konto?</strong>
 <p>
Klicka på Mitt konto och sedan på knappen Insättning i kolumnen till vänster, därefter kan du välja önskat betalningssätt.
 </p>
 </li>

 <li> <strong>Hur lång tid tar det innan min insättning blir godkänd?</strong>
 <p>
 Vid de flesta betalningssätt godkänns din insättning direkt. Vid banköverföring kan det ta upp till 7 dagar innan den når oss, och då lägger vi in insättningen på ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto.
 </p>
 </li>

 <li>
 <strong>Vilka insättningsmetoder finns tillgängliga hos er?</strong>
 <p>
Klicka på Betalningssätt överst i menyn på valfri [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sida&nbsp; för att se alla betalningssätt som är tillgängliga för dig.
 </p>
 </li>

 <li>
 <strong>Vilka kredit-/betalkort godtar ni?</strong>
 <p>
 [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] accepterar alla Visa och MasterCard/maestro kredit- och betalkort som insättningsmetoder, men det kan finnas restriktioner för uttag från MasterCard/Maestro
 </p>
 </li>

 <li>
 <strong>strong>Tillkommer det några avgifter när jag gör en insättning på mitt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto?</strong> 
 <p>
 Vi tar inte ut några avgifter när du gör insättningar på ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto.
 </p>
 </li>

 <li>
 <strong>Finns det någon lägsta/högsta beloppsgräns för en insättning?</strong> 
 <p>
 Lägsta möjliga insättning är €10 eller motsvarande i din egen valuta och högsta möjliga insättning är €5000 per dag eller motsvarande i din egen valuta.
 </p>
 </li>

 <li>
 <strong>
 Kan jag lägga in en egen gräns för insättningar per dag, vecka eller månad?
 </strong>
 <p>
 Ja, du kan lägga in insättningsgränser per Dag, Vecka och Månad. Dessa&nbsp; kan läggas in via "Mitt konto" under fliken "Ansvarsfullt spelande". Gränserna kan ändras när som helst via samma flik.
 </p>
 </li>

 <li>
 <strong>Hur gör jag en insättning från mitt bankkonto?</strong>
 <p>
 Klicka på "Insättning" i "Mitt konto" och välj Banköverföringar. Du kan aktivera det här alternativet genom att klicka på "Insättning". Följ sedan anvisningarna på skärmen.
 </p>
 </li>

 <li>
 <strong>
 Finns det någon veckogräns för hur mycket jag kan sätta in på mitt webbsideskonto via mitt bankkort?
 </strong>
 <p>Det högsta beloppet som du kan sätta in per dag är €5000.</p>
 </li>

</ol>

<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Print</span>
 </span>
 </span>
 </span>
 </button>
</p>