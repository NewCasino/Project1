Kortinnehavarens namn