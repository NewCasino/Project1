﻿[Metadata:value(/Metadata/GammingAccount/Microgaming.Display_Name)] Kredit & Debet

