Associera inte