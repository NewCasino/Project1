﻿Var vänlig skriv in beskrivning
