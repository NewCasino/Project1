﻿Om du vill begränsa ditt spelande och trappa ned, är följande alternativ möjliga för dig att inaktivera ditt konto. Notera att alla dessa alternativ är temporära. Välj en anledning nedan för att vi ska kunna förbättra din spelupplevelse. 
