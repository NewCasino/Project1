Du har just nu enastående omsättningskrav på din bonus. Om du vill ta ut eller föra över medel från {0} kontot kommer du förlora bonus eller vinster. 