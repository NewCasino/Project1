Ditt ID-nummer har redan registrerats.