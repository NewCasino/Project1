﻿minuter
