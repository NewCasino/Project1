﻿ogiltig mobil.
