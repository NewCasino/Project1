﻿Ansvarsfullt Spel
