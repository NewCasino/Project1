Fel e-postformat