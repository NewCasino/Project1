casino Bonus