Redigera bonusen T&Cs innehåll i CMS backend,/Content/Metadata/Documents/OddsMatrixTermsAndConditions