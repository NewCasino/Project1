Förbetalda kort