januari