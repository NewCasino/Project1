﻿Överför
