Felaktigt mobilnummer.