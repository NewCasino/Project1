Ogiltigt Neteller Account ID