Spela för att vinna