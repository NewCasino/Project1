﻿Registrera nytt bankkonto