För att registrera ett konto, klicka på den här länken: