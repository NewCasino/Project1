﻿Gör ett uttag direkt från din bank via DengiOnline
