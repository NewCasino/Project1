Vänligen ange Secure ID