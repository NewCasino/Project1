Fröken