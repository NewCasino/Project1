Att ta från kort nr.{0}