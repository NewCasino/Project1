Finansiella