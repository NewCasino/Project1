﻿Ditt mobilnummer här
