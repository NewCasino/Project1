﻿Adressfältet får inte lämnas tomt
