<p>Kära  $USERNAME$,<br /> </p><br />Detta e-postmeddelande får du för att bekräfta att ditt konto nu är inställt på att du är självutesluten under 6 hela månader.<br /><br /> Under denna period kommer du inte att kunna logga in på ditt konto. Vi kommer att meddela dig via e-post när perioden slutar.<br /><br />Tveka inte att kontakta oss om ni har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br /><br /><p>Kind Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kund Support Teamet</p>