﻿Din väns identitet har inte verifierats
