Ange din alias