Vänligen fyll i användarnman för TLNakit 