﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)], Cool off avslutats
