Betala per telefon (Österrike)