Ange mottagarens turkiska ID-nummer.