Sök spel via namn