Ni har uppdaterat er profil