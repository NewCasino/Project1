﻿Fel emailadress
