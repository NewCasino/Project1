﻿Förnamn måste innehålla minst två tecken
