Logga in på ditt befintliga konto