Öppna spel på en ny sida