﻿Bankkod