Direktdebitering