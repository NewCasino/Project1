Otydligt? klicka för att ändra