Sök