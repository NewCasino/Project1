﻿Reunion