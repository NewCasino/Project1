﻿/game/gamerules.jsp?game=jokerwild100&lang=sv