﻿Sidan hittades inte
