Betalningsmottagarens adress