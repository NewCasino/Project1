Spela Mynt (av Dotpay)