Nästa spel