﻿Hämtade poäng: {0}
Intjänade pengar: {1} {2}
Återstående poäng: {3}