﻿Texas hold 'em