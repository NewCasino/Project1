Söndag