﻿Meddelanden
