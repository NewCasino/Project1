﻿Account registration not allowed for single account linked vendors