﻿{0} sekunder