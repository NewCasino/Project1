Vänligen sätt in innehåll om oss här.