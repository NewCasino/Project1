Uttag av pengar direkt till ditt Clickandbuy-konto