﻿Lösenordet är inte giltig