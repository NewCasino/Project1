De kommande 6 månaderna