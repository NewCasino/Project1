Uppdatera profil