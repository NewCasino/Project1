﻿FPP Kurs
