E-postadressen matchar inte