﻿Inloggningen misslyckades. Ditt konto är under cooloff som expirerar den {0}, vänligen försök logga in då.

