Felaktigt telefonnummer.