﻿Mängd 
