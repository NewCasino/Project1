﻿/game/gamerules.jsp?game=lrcstud2&lang=sv