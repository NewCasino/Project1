﻿Populär