﻿Sätt en förlustgräns
