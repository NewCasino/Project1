Registrera med EntroPay