En 6-månaders självuteslutningsperiod