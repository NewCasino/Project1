﻿Logga ut

