<p>Hej $FIRSTNAME$,</p><p> Ditt uttag återtagits tillbaka på ‘$TXCOMPLETEDDATE$", och medlen återförts till ditt spelkonto. Kontakta support om du behöver mer hjälp angående denna transaktion.</p>Transaction ID: $TXID$Transaction Date: $TXCREATEDDATE$ Summa: $TXAMOUNT$ $TXCURRENCY$.<p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>