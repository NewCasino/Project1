Toppvinnare