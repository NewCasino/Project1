Sätt lsöenord