﻿Summa

