Avsändarens telefonnummer