﻿/game/gamerules.jsp?game=allamerican100&lang=sv