Har du frågor gällande din insättning, kontakta kundtjänsten och ange transaktions-ID-numret.