﻿Bulgariska lev
