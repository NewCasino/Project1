﻿Aktuell FPP: {0} poäng
Ｍin. poäng som krävs: {1} poäng 
Varje {2} poäng kommer att hämtas som {3} {4}

Hämta dina pengar?