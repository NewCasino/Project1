﻿Ladda ner App
