Registrera ett kort