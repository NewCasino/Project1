﻿Gått ut
