Den här kategorin innehåller dina favoritspel.