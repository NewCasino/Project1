﻿Period