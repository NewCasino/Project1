﻿Min.