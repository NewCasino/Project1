﻿Gå med nu!
