Uttagstransaktionerna som listas nedan är pågående.
Du kan ångra dessa transaktioner och återföra pengarna till ditt konto direkt genom att rycka på knappen Rulla tillbaka.
Dina pengar blir omedelbart tillgängliga på ditt konto.