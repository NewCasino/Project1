﻿Vänligen ange ditt lösenord
