Penningbelöningar