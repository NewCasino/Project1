Het