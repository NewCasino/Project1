falsk