Alla