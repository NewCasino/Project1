nummer