Ladda fler spel i den här kategorin