﻿/game/gamerules.jsp?game=victorious&lang=sv