Visa de nyaste spelen