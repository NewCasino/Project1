﻿Spela LIVE BlackJack nu!