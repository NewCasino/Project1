﻿Vänligen uppge ditt lands telefon prefix: