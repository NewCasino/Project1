Uttag direkt till ditt VISA debit kort.