<p>Kära $USERNAME$, <br /><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Syftet med detta e-mail är att bekräfta att du har ändrat din personliga förlustgräns från $LIMITAMOUNT$ $LIMITPERIOD$ till $NEWLIMITAMOUNT$ $NEWLIMITPERIOD$. <br /><br /> Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p> </p><p>Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>