Beviljat datum