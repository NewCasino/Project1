﻿/game/gamerules.jsp?game=mythicmaiden&lang=sv