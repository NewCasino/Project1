Registrera nytt bankkonto