Spelnamn