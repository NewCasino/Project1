﻿Gröntub
