Visa endast  nya bord