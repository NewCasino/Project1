Uttag direkt till ditt BOLETO konto