﻿Du har mindre än {0} i “huvudkontot”, vänligen överför tillräckligt med pengar.
