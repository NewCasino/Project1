﻿Cool-off till
