Kampanjkod