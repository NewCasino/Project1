Bekräfta