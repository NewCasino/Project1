Logga in manuellt på din internetbank och för över pengarna