Rutnät