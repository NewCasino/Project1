Vänligen ange ditt efternamn