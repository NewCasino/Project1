﻿Ta ut direkt till ditt UseMyServices konto
