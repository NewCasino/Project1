Visa alla jackpottar