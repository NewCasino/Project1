﻿Du spelar nu i {0}.