Fyll i tecknen i bilden ovan