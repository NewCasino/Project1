﻿An error has occured. Please try again later or contact support