Spelare