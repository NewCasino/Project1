Mottagarens TC nummer