Ditt förnamn innehåller ogiltiga tecken