﻿Skicka ny verifieringskod

