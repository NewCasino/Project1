﻿Möjligheter för utbetalning
