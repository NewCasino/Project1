Formatet i detta fält är ogiltigt.