﻿Bidrag till bonusomsättningen
