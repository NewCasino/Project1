﻿Transaktion historik