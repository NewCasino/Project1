Transaktionen slutförd.