spel i dina Favoriter