﻿Fyll i filialkod