﻿Fyll i ett giltigt datum 
