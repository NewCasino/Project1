﻿A technical error occurred. Invalid Mode. Please contact the merchant's customer service.