﻿Spelindex