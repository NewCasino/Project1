﻿/game/gamerules.jsp?game=arabian&lang=sv