Uttag direkt till ditt eKonto konto