﻿Blackjack US