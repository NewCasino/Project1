﻿Blackjack