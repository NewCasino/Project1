Välj det land där du är stadigvarande bosatt