Till