Vänligen ange det gamla lösenordet