Vänligen fyll i din e-post adress