Försök att utföra otillåten handling. 