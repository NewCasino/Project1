﻿ mgs-live-multispelare-blackjack
