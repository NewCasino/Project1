Ange ditt konto-ID eller din e-postadress.