Visa filter för alla kategorier