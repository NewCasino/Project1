Se alla öppningsmetoder