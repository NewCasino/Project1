Akbank är en Turkisk-baserad bank