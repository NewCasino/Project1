﻿PaymentInside