Lösenordet matchar inte