﻿Fyll i SWIFT