﻿Bordsspel

