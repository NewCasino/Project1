lägg till några spel från aktuell tillverkare.