﻿/game/gamerules.jsp?game=deuceswild10&lang=sv