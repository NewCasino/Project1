Mobilnumret matchar inte