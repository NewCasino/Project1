﻿Användarnamn:


