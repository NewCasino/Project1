﻿/game/gamerules.jsp?game=jokerwild1&lang=sv