Vi har gjort större förändringar i <a href="[Metadata:value(/Metadata/Settings.Terms_Conditions_Url)]" >Terms & Conditions</a> nyligen. Du behöver acceptera dem innan du kan fortsätta spela på vår site. Om du har några frågor vänligen kontakta vår support. 