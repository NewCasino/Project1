﻿Dölj gårdagens toppengaspelare
