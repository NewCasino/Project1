Fru