Slutdatum