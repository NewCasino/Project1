﻿För tillfället finns inga aktiva bonusar