Ogilltigt födelsedatum