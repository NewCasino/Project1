Tekniska frågor