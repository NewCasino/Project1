Uppdatera