﻿Verifieringskoden misslyckades att skickas, kontrollera ditt telefonnummer eller försök igen.

