﻿/game/gamerules.jsp?game=cstud2&lang=sv