Öppna spel på den här sidan