﻿Konto-ID/E-postadress