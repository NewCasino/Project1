Vänligen ange ditt konto ID