Spelegenskaper: