﻿Neteller(Bulgarien)
