Tyvärr, länken är för gammal eller ogiltig.