E-postmeddelandet kunde inte skickas just nu. Försök igen senare.