Uttag av pengar direkt till ditt Poli-konto