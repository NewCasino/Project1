﻿Glömt Lösenord
