﻿Klassiska automater
