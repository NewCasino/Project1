﻿Lista