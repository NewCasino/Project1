﻿Registrera  ett kort
