E-plånböcker