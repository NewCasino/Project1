Ansvarsfullt spelande