Avvisa