﻿Självexkludera till
