Ange din kompis e-postadress.