﻿Uttag från