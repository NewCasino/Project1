TILLGÄNGLIGA BONUSAR