Tisdag