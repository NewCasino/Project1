﻿Reklamerade Poäng: {0}<br/>Tjönade Pengar: {1} {2}<br/>Återstående punkter: {3}
