Lär dig mer om belöningar