Spela på skoj