﻿/game/gamerules.jsp?game=blackjackdblex&lang=sv