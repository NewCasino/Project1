﻿För din säkerhet ber vi dig ändra ditt lösenord för att följa de nya lösenordsreglerna.
