﻿Tidszon
