﻿Lägga till {0}  hemskärm
