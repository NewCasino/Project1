﻿OBS! Du får bara växla in <span class='messageHighlight'>{0}</span> poäng för 
<span class='messageHighlight'>{1} {2}</span>. Återstående poäng kommer att stanna kvar på ditt FPP-konto.

