Du hamnade troligen på den här sidan av misstag.