<p>$FIRSTNAME$,</p><p> Para yatırma talebiniz başarısız olmuştur. Lütfen bilglierinizi kontrol edip tekrar talep verin.</p><p> Lütfen herhangi bir problem yaşadığınız taktirde aşağıdaki email adresinden müşteri hizmetlerine başvurunuz: </p><p><a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a> .<br /> <br /> Saygılarımızla ,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]</p>