﻿Ditt postnummer här
