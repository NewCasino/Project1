﻿Vi beklagar men du är inte berättigad att göra en överföring just nu. Vänligen <a href="/ContactUs">kontakta kundtjänst</a> för ytterligare information.