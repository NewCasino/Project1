﻿/game/gamerules.jsp?game=reelpoker&lang=sv