månad