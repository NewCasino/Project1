﻿Välj bonus
