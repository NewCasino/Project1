﻿Smart SMS-lösenord