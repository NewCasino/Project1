<p> Hi $FIRSTNAME$, </p> Din utbetalning för $VOUCHERAMOUNT$ har bearbetats. Nedan finns information om din IPS Token:</p><ul><li><strong>IPS Token</strong>:$VOUCHERNUMBER$</li><li><strong>Checkdigit</strong>:$VOUCHEDIGITS$</li></ul><p>Om du har några frågor tveka inte att kontakta<a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Vänligen,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>