﻿Nedtrappning under 7 dagar
