﻿/game/gamerules.jsp?game=allamerican10&lang=sv