﻿Kasino Information
