﻿Yandex.Money är ett betalningssystem som tillåter deras användare att betala och ta emot betalningar online via webb samspel, smarttelefoner och tablettapplicationer.
