﻿/game/gamerules.jsp?game=retro-super80&lang=sv