Captcha är inkorrekt, vänligen försök igen. 