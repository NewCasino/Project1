Med ﻿POLi by Skrill kan du föra över pengar från en bank direkt till ditt konto. Du behöver inte vänta på att pengarna ska klareras, betalningen sker direkt.&nbsp;POLi är ett av Australiens effektivaste betalningssätten online.