﻿Dubbel Bonus Serier
