﻿Uttag till ett annat konto
