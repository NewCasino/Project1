﻿Användar-ID
