﻿Inträde
