﻿Frankenstein™ är ett 5 reel, 3 rad och 20 bet line video slot med maxsatsning på € 100. Det intruduserar nya utseendetLinked Wilds™som framträder i båda huvudspelen och Free Spinns.
