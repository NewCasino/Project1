Välj en tillverkare: