E-postadressen är inte tillgänglig eller har redan tagits av någon annan, försök med en annan e-postadress.