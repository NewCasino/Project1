﻿Banköverföring

