﻿Text:
