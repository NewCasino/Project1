﻿Sätt en omsättningsgräns
