Dealerns ursprung