﻿Profil