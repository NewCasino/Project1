﻿Casinospel - Bonuspremie