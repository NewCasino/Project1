Ändra maxbelopp