Jag har läst och bekräftat meddelandet ovan.