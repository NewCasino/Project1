﻿Jacks eller Better Serier

