Hem