Ange ditt gamla lösenord