﻿Välj Kreditkort
