﻿Bonuskontrib.
