<p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] har förbundit sig att stödja ansvarsfullt spelande som ett sätt till kundvård och socialt ansvar. Vi tror att det är vårt ansvar gentemot dig, våra kunder, att se till att du njuter av din spelupplevelse på vår webbplats. <br /> <br />Spel bör ses som ett roligt tidsfördriv, och inte som ett sätt att generera intäkter. Medan majoriteten av befolkningen kan behandla spelandet som rekreation och spenderar bara vad de har råd att riskera, kan det för vissa vara svårare. För att upprätthålla kontrollen över dina spelvanor vill vi påminna dig om att alltid tänka på följande punkter:  <br /> <br />* Spelande bör göras med måtta och genomförs som en form av fritid inte som ett äkta sätt att tjäna pengar <br />* Undvik att jaga förluster - det kommer alltid att komma en ny dag.<br />* Spela endast så du kan täcka förlusterna <br />* Håll koll på tiden och övervaka mängden pengar du spenderar <br />* Skulle du behöva en paus från spelandet, kan själv-uteslutning från ett eller alla produkter aktiveras genom att kontakta Support. <br /> <br />Om du behöver prata med någon om eventuella problem du kan ha med ditt spelande, vänligen kontakta någon av de organisationer som vi har listat nedan.</p><br /><p><strong>Har du ett problem ?</strong> <br /> <br />Om du är orolig för att spelandet har haft en negativ inverkan på ditt eller någon annans liv kan följande frågor hjälpa dig. <br /> <br />1. Hindrar spelet dig från att gå jobbet eller skolan <br />2. Spelar du för att fördriva tiden eller att fly tristess? <br />3. Spelar du ensam under långa perioder? <br />4. Har andra kritiserat någonsin dig för ditt spelande? <br />5. Har du förlorat intresset för familjen, vänner eller fritidsintressen pga spelande? <br />6. Har du någonsin ljugit för att dölja hur mycket pengar eller tid du spenderar på spelandet? <br />7.Har du ljugit, stulit eller lånat för att upprätthålla dina vadslagnings vanor? <br />8. Är du tveksam till att spendera "spelpengar" på något annat? <br />9. Spelar du tills du förlorar alla dina pengar? <br />10. Efter att ha förlorat, känner du att du måste försöka vinna tillbaka förlusterna så fort som möjligt? <br />11.Om du får slut på pengar när du spelar, känner du dig vilsen och förtvivlad och känner behov av att spela igen så snart som möjligt? <br />12. Gör gräl, frustration eller besvikelser att du vill spela? <br />13. Gör spelande dig deprimerad eller självmordsbenägen? <br /> <br />Ju fler frågor som du svarar "ja" till, desto mer sannolikt är det att du har problem med ditt spelande. Att prata med någon som kan ge dig råd och stöd, vänligen kontakta någon av de organisationer som anges nedan under Organisationer Gambling Rådgivning.</p><br /><p><strong>Insättningsgränser</strong> <br /> <br />för att hjälpa våra spelare i spel på ett ansvarsfullt sätt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] finns det en insättningsgräns möjlig på varje kundkonto. Denna möjlighet finns tillgänglig under "<a href="/profile">My Account</a>". Gränser kan ändras när som helst. En minskning av depositionsgränsen träder i kraft omedelbart, men en ökning kan endast ske efter en betänketid, för att undvika förhastade beslut.<br /> <br />Om du behöver ytterligare information eller hjälp gällande  funktionen, kontakta <a href="/contactus">Support</a>.</p><br /><p><strong>Self-exclusion</strong> <br /> <br />Om du behöver ta en paus från spelandet, tillhandahåller vi en<a href="/SelfExclusion">självuteslutning</a>åtgärd som kan aktiveras av kunden under "Mitt konto" eller genom att kontakta support. Självuteslutning innebär att ditt konto kommer förbli stängt under en period av minst 7 dagar, och kommer inte att återaktiveras under några omständigheter under uteslutningsperioden. Detta är den stora skillnaden för när du avslutar ett konto på "vanligt" sätt. En skriftlig begäran (upphör efter din angivna tidsramen) krävs innan kontot återöppnande kan övervägas. <br /> <br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]  ger kunderna möjlighet att blockera åtkomst till enskilda produkter (Sportsbook, Casino Games och Poker) via "Mitt konto" eller genom att kontakta support  <br /> <br />Om du funderar självuteslutning, kom ihåg att kontakta alla spelbolag som du har konton och begära att självuteslutning hos dem också. Vi rekommenderar också att du tänker på en eventuell installation av programvara som gör att du kan blockera åtkomst till webbplatser. Se filtreringssystem längst ner på denna sida. </p><br /><p><strong>Gambling Counselling Organisations</strong> <br /> <br />* GamCare, den ledande auktoriteten för att erbjuda rådgivning och praktisk hjälp i hanteringen av sociala effekterna av spelande i Storbritannien, kan besökas på: www.gamcare.org.uk . Dess konfidentiella hjälplinje är: 0845 6000 133. Icke - brittiska medborgare kan kontakta GamCare för information om internationella stödorganisationer. <br />* Gamblers Anonymous är en gemenskap av män och kvinnor som har gått samman för att göra något åt ​​sina egna spelproblem och hjälpa andra spelmissbrukare att göra detsamma. Det finns regionala stipendier runt om i världe . Gamblers Anonymous internationella tjänst webbplats är: www.gamblersanonymous.org.uk. </p><br /><p><strong>Minderåriga spel</strong> <br /> <br />Det är olagligt för någon under 18 år att öppna konto och spela på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]  tar sitt ansvar gällande detta mycket allvarligt och förutom våra slumpvisa kontroller gällande ålder, genomgör vi åldersverifikation på alla spelare som använder betalningsmetoder som användar eunder 18 år kan göra. Vi förbehåller oss rätter att fråga efter dokumentation som kan verifiera din ålder, och ditt konto kommer att stängas av fram till att dokumentation kan uppvisas </p><p> </p><p>Om du delar dator med vänner eller familj som är under 18 rekommenderar vi lösningar så som filter för föräldrakontroll, sådan programvara tillåter föräldrar att reglera tillgång till Internet för att barn inte ska kunna ha tillgång till spelsidor online. </p><p> </p><p>Net Nanny™ www.netnanny.com</p><p>CyberPatrol www.cyberpatrol.com</p><button type="button" onclick="window.print(); return false" class="button"> <span class="button_Right"> <span class="button_Left"> <span class="button_Center"> <span>Print</span> </span> </span> </span> </button></p>