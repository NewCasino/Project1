Veckogräns (per vecka)