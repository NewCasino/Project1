﻿/game/gamerules.jsp?game=robinhood&lang=sv