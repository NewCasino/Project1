﻿/game/gamerules.jsp?game=tiki&lang=sv