﻿Välkommen till 

