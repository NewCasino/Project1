Villkor