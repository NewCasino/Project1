Månatlig gräns (per månad)