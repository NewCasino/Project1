Byt lösenord