De kommande 7 dagarna