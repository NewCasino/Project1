Vänligen ange ett nytt lösenord