﻿/game/gamerules.jsp?game=lrblackjackmini&lang=sv