Inloggningen misslyckades. Ditt användarkonto är blockerat.
Om du är en självutesluten användare, kontakta kundtjänst för hjälp med uttag av pengar