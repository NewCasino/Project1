﻿/game/gamerules.jsp?game=fruitshop&lang=sv