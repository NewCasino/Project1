Login misslyckades. Ditt konto är blockad.Om du har självblockad dig kontot, vänligen kontakta supporten