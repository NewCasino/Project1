﻿Ange bonuskod
