Ange verifieringskod