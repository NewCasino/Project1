<p>$FIRSTNAME$,</p><p> Para yatırma talebiniz onaylanmıştır, [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] 'i seçtiğiniz için teşekkür eder, oyunlarımızda bol şans dileriz. </p><p> Lütfen herhangi bir problem yaşadığınız taktirde aşağıdaki email adresinden müşteri hizmetlerine başvurunuz:</p><p> <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a> .</p><p> Saygılarımızla ,</p><p> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]</p>