Affiliate-markören kommer att trunkeras eftersom dess längd överstiger gränsen.