Ditt land stöds inte, försök använda andra metoder