﻿Du har redan loggat in [Metadata:value(/Metadata/Settings.Operator_DisplayName)].