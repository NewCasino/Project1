﻿Observera att meddelandenumret bara kan endast användas vid en insättning. Den andra insättningen med samma meddelandenummer kommer inte att fungera.

