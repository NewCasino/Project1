Verifkationstext ogiltig, försök igen