Bekräfta e-postadressen