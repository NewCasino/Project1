﻿Starta