﻿Bearbetar

