﻿Överföring till användar- {0} {1} konto