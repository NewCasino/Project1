Spela