﻿Belopp
