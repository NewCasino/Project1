﻿Du går in på mobila upplagan, vill du byta till Skrivbord Edition?
