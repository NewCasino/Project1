﻿/game/gamerules.jsp?game=tfhvideopokerdw&lang=sv