Visa spel i rutnätsvy