Användarmeddelanden 