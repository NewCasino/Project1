Endast män