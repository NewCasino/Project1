Nytt lösenord