﻿Användarnamnet måste väljas
