﻿Vänligen ange ditt citizen ID
