Bank of Georgia (bankomat)