﻿Fisticuffs
