﻿All American Serier
