Lägg in spelets namn: