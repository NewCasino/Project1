﻿Namn på konto
