﻿Cancellation declined - no reference ID.