Du måste logga in för att genomföra aktiviteten.