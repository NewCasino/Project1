﻿Vänligen välj en vän att överföra till.
