Spela på låtsas