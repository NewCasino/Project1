Du måste bekräfta att du accepterar våra villkor och bestämmelser