﻿Buddy transfer