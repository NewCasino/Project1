Fel lösenord.