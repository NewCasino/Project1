﻿Transaktionen ej tillåten!
