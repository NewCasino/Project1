﻿falsk