﻿Neteller(Denmark)