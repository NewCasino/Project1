﻿Sportsbooks Regler