﻿Oddsformat
