﻿/game/gamerules.jsp?game=blackjackonedk&lang=sv