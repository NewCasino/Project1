﻿Överföring av pengar direkt till ditt bankkonto

