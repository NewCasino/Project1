﻿/game/gamerules.jsp?game=hrhilo&lang=sv