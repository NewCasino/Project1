﻿Vunna spel
