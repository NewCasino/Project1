Ukash nummer