Din förfrågan att återställa detta uttag kan inte bearbetas för tillfället. 