﻿<ol>

 <li> <strong>Hur kan jag identifiera betalningar eller uttag till [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] på mitt bank/kreditkortsutdrag?</strong> 
 <p>
 Alla insättningar och uttag&nbsp; på ditt kredit- eller bankkontoutdrag visas tillsammans med en deskriptor där [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] anges. Det gör att du kan hålla koll på dina insättningar till och uttag från sidan.
 </p>
 </li>

 <li> <strKan jag använda mer än ett betalningssätt?</strong>
 <p>*Ja, det kan du, men vi kan behöva dokumentation vid ändring av betalningssätt.
 </p>
 </li>

 <li>
 <strong>Accepterar ni kort från mitt land?</strong>
 <p>*Vi accepterar kort från alla länder utom USA, Turkiet och Frankrike.
 </p>
 </li>

 <li>
 <strong>Varför acceptera er webbsida inte mitt kort?</strong>
 <p>
Vissa kreditkortsutgivare har som regel att inte tillåta direktbetalningar till spelsidor online. Du kan kontakta din kortutgivare angående detta eller försöka göra en insättning via en e-plånbok istället.&nbsp; För ytterliga hjälp kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kundtjänst.
 </p>
 </li>

 <li>
 <strong>Vad gör jag om min kortinsättning inte accepteras eller avslås?</strong>
 <p>
Om du försöker göra en andra insättning bara en kort stund efter det att en föregående insättning gått igenom kan det hända att den räknas in i din 24-timmars eller veckovisa insättningsgräns, vilket orsakar insättningsproblem. Den vanligaste orsaken till att problemet uppstår är dock att fälten i ansökningsformuläret inte har fyllts i korrekt. Kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kundtjänst för att rätta till problemet. Vissa kreditkortsutgivare har också som regel att inte tillåta direktbetalningar till spelsidor online. Du kan kontakta din kortutgivare angående detta eller försöka göra en insättning via en e-plånbok istället.
 </p>
 </li>

 <li>
 <strong>Kan jag använda mitt kort för att göra en insättning på en kompis konto?</strong>
 <p>
Det kan du inte göra eftersom det anses som en tredjeparts-transaktion och är under inga omständigheter tillåtet.
 </p>
 </li>

 <li>
 <strong>Jag har av misstag satt in pengar från fel kort &ndash; vad gör jag?</strong> 
 <p>
Kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst
 <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">
 [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]
 </a>
 </p>
 </li>

 <li>
 <strong>Kan jag föra över pengar mellan konton?</strong>
 <p>
Du kan inte föra över pengar mellan personliga konton men du kan föra över pengar mellan Casino, Sports Book och Poker i ditt personliga konto.
 </p>
 </li>

 <li>
 <strong>Vad är en IBAN?</strong>
 <p>
IBAN står för International Bank Account Number. IBAN används vid internationella banköverföringar och gör det enklare för dig att ta ut dina vinster.
 </p>
 </li>

 <li>
 <strong>Vad är en CVC2?</strong>
 <p>
CVC2 är en akronym för "Card Verification Code". Den här koden krävs som en säkerhetsåtgärd när du gör internationella telefonköp och internetbetalningar med bankkort. Den här koden består av tre siffror och finns på baksidan av ditt bankkort.
 </p>
 </li>

</ol>

<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Skriv ut</span>
 </span>
 </span>
 </span>
 </button>
</p>