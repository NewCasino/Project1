﻿Visa Balansen
