﻿Vänligen skriv in din väns E-post
