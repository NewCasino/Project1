﻿Inloggning lyckades. Du kommer inom kort omdirigeras.
