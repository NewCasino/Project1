Belopp som ska föras över till {0}