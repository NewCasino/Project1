﻿/game/gamerules.jsp?game=hrtreypoker-1h&lang=sv