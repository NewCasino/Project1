﻿Säkert
