﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Ditt uttags IPS-kvittens