Alla vinnare