﻿Saldo
