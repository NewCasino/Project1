Du kommer inte kunna logga in på ditt vadslagningskonto under en period av 3 månaders avkylning.