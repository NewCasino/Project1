﻿Vänligen bekräfta ditt lösenord
