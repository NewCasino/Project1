Tekniska problem