﻿Säkerhetskod
