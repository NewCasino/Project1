Uttag av pengar direkt till ditt Click2Pay-konto