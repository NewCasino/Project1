Fel uppstod.