juni