Kära $USERNAME$, <br /><br /> Syftet med detta e-mailet är till för att bekräfta att perioden av ditt permanenta självutslutnings period nu har avslutas och att alla funktioner på ditt konto nu är tillgängliga. <br /><br />Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Vänliga hälsningar </p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Customer Support Team</p>