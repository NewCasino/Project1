﻿<ul>
<li>
<strong>Privat Policy</strong>
<p>
Genom att använda och eller besöka några sektoner på webbsidan [Metadata:value(/Metadata/Settings.Operator_DisplayName)] (the <b>"Website"</b>); eller öppna ett konto på webbsidan godkänner du den privata policyn. Vid användning av webbsidans produkter kommer du att blitillfrågan att överlämna oss med riktig, uppdaterad personuppgifter som kommer tllåta oss att identifiera dig.</p>

<p>
i) Du implicit ge ditt tillstånd till behandling av personuppgifter i enlighet med sekretesslagar i tillämliga jurisdiktioner.</p>
<p>
ii) Du bekräftar din vilja att dela med dig av särskild privat information me företaget som kommer att används för att bekräfta din identitet. Denna information samlas i linje med våra stränga kontrollförfaranden som används för att avskräcka internationella penningtvätt och för att säkerställa säkerheten för spelarnas aktivitet.</p>
<p>
Företaget har åtagit sig att skydda och respektera din integritet, sekretessoch säkerhet och att fullt ut följa dataskydd och sekretesslagar. </p>
</li>
<li>
<strong>Samling av Personuppgifter: </strong>
<p>Vi samlar in denna information när du registrerar dig och använda våra spelprodukter, göra förfrågningar, anmälsa sig till erbjudanden eller andra tjänster eller när du besvarar kommunikation från oss såom, men inte begränsat till undersökningr och frågor
. Den information vi samlar in kan inkludera personlig och bankuppgifter och all annan information som du delar dig med oss.</p> 
</li>
<li>
<strong>Hur denna information behandlas</strong>
<p>Den information
 du ger oss kommer att behandlas för ett antal skäl, däribland att tillhandahålla dig med peltjänster, för att behandla ansökningar du gör för informatio för att förse dig med tillräckligt stöd, av marknadsföringsskäl, att meddela dig om eventuella ändringar vi kan göra vår tjänst eller webbplats från tid till en annan för att uppfylla de skyldigheter som åläggs av tillsynsmyndigehter i jurisdiktioner där vi har e licens och för någon av de speciferade anledningen till att du ombads att lämna uppgifter om. </p>
</li>
<li>
<strong>Vilka lämnar vi ut din personuppgifter till: </strong>
<p>
Dina personuppgifter kan lämnas ut till:<br />
a)  Bolag inom koncernen. I detta fall ser vi till att endast behöriga anställda får tillgåg till det;<br />
b) Till tredjepartsföretagen som driver ett white label varumärke med hjälp av våra tjänster och ge dig speltjänster;<br />
c)  Till tredjeparts företagsom tillhandahåller tjänstertill vårt företag som i sin tur hjälper oss att leverera speltjänster, men inte begränsat till betalning processorer eller datakontrollanter;<br />
d)  Till konsulter såsom reisorer som erbjuder sina tjänster till företag eller något företag inom vår gruppoch som är avsedda att hjälpa os att bättra vår verksamhet;<br />
e)  Till eventuella investerare eller köpare av alla företag som ingår i koncernen;<br />
f)  Till statliga myndigheter eller insitutioner men denna överföring kommer skekrävs  endast med särskild med lagen.<br />Någon tredje part som vi väljer att avslöja dina personuppgifter till kommer att vara avtals skyldiga att följa dataskydd och integritetslagar och villkoren i denna integritetspolicy
. </p>
</li>
<li>
<strong>Säkerhet</strong>
<p>Företaget lovar att vidta åtgärder och politik som hjälper till att skydda din personliga information från obehörig åtkomst eller obehöriga ändringar, avslöjanden eller förstörelse
.</p>

<p>
Du kan skriva till oss på <a href="mailto:[Metadata:value(/Metadata/Settings.Email_SupportAddress)]">[Metadata:value(/Metadata/Settings.Email_SupportAddress)]</a>  om du vill få en kopi av dina personuppgifer eller om du vill ändra dina personuppgifter på något vis.</p>
</li>
<li>
<strong>Miscellaneous</strong>
<p>
Dina personuppgifter kommer att hållas av oss så länge som det tjänar syftet till att densamlades in.</p>

<p>
Vi har rätten att modifiera eller ändra denna integritetspolicy då och då. I den ossannolika händelse av ändringar görs kommer vi att meddela dig så nart som möjligt och vid behov kommer vi att fråga om ditt samtycke.</p>

<p>
Om du har några funderingar kring vår privatpolicy, vänligen skriv till oss på <a href="mailto:[Metadata:value(/Metadata/Settings.Email_SupportAddress)]">[Metadata:value(/Metadata/Settings.Email_SupportAddress)]</a>.</p>
</li>
</ul>
<p style="text-align: right">
    <button class="button button-print" onclick="window.print(); return false" type="button">
        <span class="button_Right"><span class="button_Left"><span class="button_Center"><span>
            Print</span> </span></span></span>
    </button>
</p>




