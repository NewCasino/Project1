Du har blivit frånkopplad då någon har loggat in med ditt konto på en annan plats. Var vänligen notera att om detta inte var avsiktligt kan någon ha stulit ditt lösenord och vi föreslår att du ändrar det omedelbart.