<p>Kära $USERNAME$,<br /></p><br />Syftet med detta e-mail är att bekräfta att ditt konto nu är inställd på självutslutning under perioden av 1 år.<br /><br />Under den här perioden kommer du inte kunna logga in på ditt konto. Vi kommer meddela dig via e-mail när perioden av självutslutning är över.<br /><br />Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br /><br /><p>Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>