Uttag direkt till ditt Maestro kort.