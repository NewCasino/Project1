﻿Referens