Snabb banköverföring