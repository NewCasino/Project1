Växlingssumma: