Lösenordet saknas