Välj giltighetstid t.o.m.