﻿Japan, Japanese Yen