Observera att gränserna är baserade på kalendervecka eller -månad. Angivna insättningsgränser återställs i början av varje vecka eller månad. Exempel: Om du har angett en insättningsgräns på € 100 den 20 augusti och sätter in maxbeloppet i slutet av månaden, kan du sätta in € 100 igen fr.o.m. den 1 september.