﻿Vouchernummer krävs
