Uttag direkt till ditt Click2Pay konto