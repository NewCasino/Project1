﻿Ogiltigt UIPAS Konto ID.
