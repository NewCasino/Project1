Uttag direkt till ditt GiroPay konto