﻿Bettinghistorik
