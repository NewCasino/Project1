Se alla jackpottar nu!