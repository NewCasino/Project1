﻿Valideringskoden krävs
