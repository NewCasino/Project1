Spela nu!