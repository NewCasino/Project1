﻿Ange token
