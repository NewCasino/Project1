Beloppet kan inte vara tomt.