Bankkontonumret används redan, välj ett annat