﻿Bekräftelse
