﻿Alla Americans II
