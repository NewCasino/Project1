﻿<ol>

    <li> <strong>Var är er webbsida baserad?</strong>
        <p>Vår webbsida är baserad på Malta.</p>
    </li>

    <li> <strong>Är er webbsida licensierad?</strong>
        <p>
            Ja, vi har en giltig EU-licens för spel på sport, casino och poker.
        </p>
    </li>

    <li>
        <strong>Hur säkra är mina bankkortsuppgifter?</strong>
        <p>
            [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] använder de mest avancerade kryperingsteknikerna för att garantera att dina uppgifter endast är tillgängliga för några få utvalda inom [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] familjen. Vi krypterar alla dina uppgifter med hjälp av krypteringsalgoritmer enligt den internationellt godkända standarden SSL. Det gäller alla dina uppgifter som skickas fram och tillbaka; från din adress, till korten som du tilldelats hanteras med lika hög skyddsnivå som en bank skulle använda.
        </p>
    </li>

    <li>
        <strong>Hur vet jag att mina finansiella uppgifter är säkra?</strong>
        <p>
            [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] krypterar alla dina uppgifter med hjälp av krypteringsalgoritmer enligt den internationellt godkända standarden SSL. Det gäller alla dina uppgifter som går fram och tillbaka; från din adress, till korten som du tilldelats hanteras med samma skyddsnivå som den säkerhet som en bank använder.
        </p>
    </li>

    <li>
        <strong>Hur vet jag att mina pengar är säkra?</strong>
        <p>
            Alla kundmedel sätts in på ett separat kundmedelskonto på Bank of Valetta. Detta sker i enlighet med Maltas bestämmelser för lotterier och spel, där vi även är licensierade. Kundmedlen hålls helt "isolerade" från företagets medel och förvaras säkert på det här sättet för att säkerställa att kundmedlen alltid finns tillgängliga för våra kunder.
        </p>
    </li>

</ol>

<p style="text-align:right">
    <button type="button" onclick="window.print(); return false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span>Print</span>
                </span>
            </span>
        </span>
    </button>
</p>