Uttag direkt till ditt eWire konto