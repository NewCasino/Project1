﻿Neteller(Ukraina)
