Är du säker på att du vill ta bort gränsen?