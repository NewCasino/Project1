Ange ditt konto-ID/din e-postadress