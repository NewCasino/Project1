Sök spel...