﻿Casino-bonus