﻿Videospelautomater
