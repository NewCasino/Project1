﻿Bonus erbjudande
