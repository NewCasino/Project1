TLNakit användarnamn