﻿Du har loggatsut automatiskt för du har varit inaktiv förlänge. Av säkerhetsskäl har du blivit utloggad automatiskt. Vänligen klicka OK för att logga in igen
.

