﻿Ta ut direkt till din bank med Alternative Payment Exchange
