﻿Välj ett spelkonto.
