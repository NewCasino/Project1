﻿/game/gamerules.jsp?game=lostpyramid&lang=sv