Min favoirtfärg?