﻿/game/gamerules.jsp?game=lrpuntobanco&lang=sv