Lösenordet måste bestå av bokstäver och siffror.