﻿Inbetalning med
