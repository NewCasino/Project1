Vänligen välj vilket datum giltigt till.