﻿Adress linje 1
