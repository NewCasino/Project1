﻿Postnummer måste anges
