Inloggningen misslyckades. Du har inte aktiverat ditt konto.