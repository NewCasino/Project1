Ange plånbokens nummer.