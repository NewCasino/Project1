﻿/game/gamerules.jsp?game=excalibur&lang=sv