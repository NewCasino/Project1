﻿Härmed bekräftar jag att jag är 18 år eller äldre och godkänner regler och villkor
