﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Bytningen av Ukash kupong
