Favoriter