﻿/game/gamerules.jsp?game=shoot4gold&lang=sv