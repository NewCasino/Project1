﻿Demospel
