﻿Konto holding filial