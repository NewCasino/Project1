Du har blivit frånkopplad då din begränsade sittningstid har nåtts.