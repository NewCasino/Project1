Klicka för att spela