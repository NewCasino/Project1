schweizisk Franc