Gör ett uttag direkt till ditt WebMoney konto