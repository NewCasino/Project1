﻿spel/sida