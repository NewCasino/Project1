﻿Lösenordet får inte vara det samma som användarnamnet.
