Slumpmässigt bord