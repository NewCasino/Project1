﻿Zimpler