Ange betalningsmottagarens adress.