Repeterade lösenordet fattas