﻿Efternamn
