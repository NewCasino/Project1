Betala per telefon (UK)