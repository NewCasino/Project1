﻿Casino poäng för frekventa spelare
