﻿/game/gamerules.jsp?game=troll&lang=sv