﻿Uttag direkt till ditt bankkonto.
