Ditt svar måste bestå av minst 2 tecken