﻿Avbryt Uttag