﻿<ol>

 <li> <strong>Har ni någon min- och maxgräns för insatser?</strong>
 <p>** Maxgränsen varierar beroende på evenemanget. Om du försöker satsa mer än maxgränsen, får du ett meddelande som talar om vilket maxbelopp du kan satsa på ditt val. Vi har ingen minimigräns för insatser.
 </p>
 </li>

 <li> <strong>Vad är enskilda insatser och multipla insatser?</strong>
 <p>
En enstaka insats gäller just ett val; en multipel insats kräver mer än ett. Ju fler val du länkar ihop i en multipel (t.ex. alla hemmalag i en omgång av Premier League), desto mer kan du vinna&ndash; men så är det ju mycket svårare!
 </p>
 </li>

 <li>
 <strong>Hur många val kan ingå i en multipel insats?</strong>
 <p>
 Det maximala antalet alternativ som vi tillåter vid multipla insatser är 10.
 </p>
 </li>

 <li>
 <strong>Hur fungera handikappbetting?</strong>
 <p>
 För detaljerad beskrivning av handicap-betting (1x2 med Handicap och Asiatiska handicap), besök avsnittet för bettingbeskrivning här.
 </p>
 </li>

 <li>
 <strong>Vad händer om en match blir uppskjuten?</strong>
 <p>
 Kontrollera reglerna för den sporten. Vissa sporter kräver att matchen spelas på samma dag för att insatsen ska bestå, insatser i andra sporter kan förbli öppna tills matchen har slutförts eller officiellt blivit stoppad.
 </p>
 </li>

 <li>
 <strong>Varför har min vinnande insats inte betalats ut ännu?</strong>
 <p>
 [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] kräver att officiella resultat har meddelats innan utdelningen kan fastställas. Ibland kan onlinekällor som live poängsajter vara felaktiga varför utdelningen kan bli fördröjd tills resultaten kan bekräftas.
 </p>
 </li>

 <li>
 <strong>Jag har ändrat mig, kan jag ångra min insats?</strong>
 <p>
 Nej, när du väl har bekräftat din insats och den har accepterats av din server, kan du inte ta tillbaka den.
 </p>
 </li>

 <li>
 <strong>Var kan jag hitta en lista över mina insatser?</strong>
 <p>
 Din insats- och transaktionshistorik finns under "Mitt sportsbetting-konto" när du är inloggad på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sajten.
 </p>
 </li>

 <li>
 <strong>Varför beräknas vinsterna annorlunda på UK-odds?</strong>
 <p>
Vid beräkningen av vinster, använder vid decimal (EU) odds eftersom de är mer exakta. UK- och US-odds är endast avsedda för visning eftersom vissa decimal-odds inte korrelerar med en enkel fraktion.
 </p>
 </li>

 <li>
 <strong>Betting börjar bli vanebildande för mig, vad gör jag?</strong>
 <p>
 Betting med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] ska vara en trevlig fritidssysselsättning för alla, men för en liten grupp människor kan det bli ett beroende och skapa problem. Information om spelmissbruk finns under Ansvarsfullt spelande.
 </p>
 </li>

</ol>
<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Print</span>
 </span>
 </span>
 </span>
 </button>
</p>