﻿<ol>
  <li><strong>Var hittar jag aktuella kampanjer?</strong>
    <p>Du hittar alla aktuella kampanjer genom att klicka på vår [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kampanjer-flik.</p>
  </li>
  <li><strong>Kan jag spela alla spel på webbsidan när jag får en bonus, eller finns det begränsningar för vilka spel jag kan spela?</strong>
    <p>Läs igenom villkor och bestämmelser för bonus och om du har frågor kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] vår kundtjänst.</p>
  </li>
  <li><strong>Hur kontrollerar jag om jag uppfyller kraven för en utdelning?</strong>
    <p>Du kan kontrollera dina framsteg genom att klicka på "mitt konto", därefter på mitt sport-konto på vänster sida och sedan på aktiva kampanjer.</p>
  </li>
  <li><strong>Varför blir jag nekad utdelning?</strong>
    <p>Vissa kampanjer gäller endast för personer från vissa länder och vissa kunder som använder specifika betalningssätt. Det kan finnas begränsningar för vissa länkade konton och missbruk av [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] utdelningar, för ytterligare anvisningar kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p>
  </li>
</ol>
<p style="text-align:right">
  <button type="button" onclick="window.print(); return false" class="button"> <span class="button_Right"> <span class="button_Left"> <span class="button_Center"> <span>Skriv ut</span> </span> </span> </span> </button>
</p>