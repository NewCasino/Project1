Skriv in kontrollsiffrorna.