En permanent självutslutningsperiod