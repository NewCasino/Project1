Ditt säkerhets-ID måste bestå av minst 6 tecken