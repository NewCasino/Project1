﻿Oddshistorik
