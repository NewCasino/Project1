[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Återställ ditt lösenord