Kort-värde