Välj en fråga