Uttag av pengar direkt till ditt bankkonto