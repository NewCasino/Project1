Beviljandedatum