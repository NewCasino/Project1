﻿Kontakta oss
