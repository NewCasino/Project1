﻿Jackpot Spel
