﻿Frankenstein™
