﻿Fruit Bonanza
