Associera