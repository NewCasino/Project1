Valuta och belopp