﻿<span class="TotalGameNumber">{0}+</span> Spel