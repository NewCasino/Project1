﻿Logga in på ditt konto


