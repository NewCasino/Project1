Du kommer inte kunna logga in på ditt konto under de nästkommande 7 dagarna