﻿Inga uppgifter kunde hittas
