﻿/game/gamerules.jsp?game=dragonisland&lang=sv