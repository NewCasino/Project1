﻿/game/gamerules.jsp?game=lrtxsholdem&lang=sv