Uttag av pengar direkt till ditt MULTIBANCO-konto