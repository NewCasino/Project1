Transaktionen har återtagits.