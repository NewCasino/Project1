Polen, Zlotych