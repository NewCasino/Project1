﻿Captcha är fel. Försök igen!

