Uttag direkt till ditt bank konto