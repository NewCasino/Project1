﻿Skraplotter
