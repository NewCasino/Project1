﻿Logga in
