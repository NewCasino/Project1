Förlustgräns