﻿Todito-kort