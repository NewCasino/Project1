﻿MULTIBANCO