Visa de populäraste spelen