Försök till icke godkänd operation.