Vänligen välj valuta