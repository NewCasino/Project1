﻿United Kingdom