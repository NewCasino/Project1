Venezuela Bolivar Fuerte