﻿Banknamn