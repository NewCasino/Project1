Stäng det här popupfönstret nu!