Vänligen ange tecknen in bilden