EWIREDK