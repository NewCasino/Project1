Dölj stängda bord