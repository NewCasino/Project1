Uttag av pengar direkt till ditt Switch/Solo-kort.