Kreditera {0} konto.