﻿[metadata:value(/Deposit/_Index_aspx.Tab_RecentPayCards)]
