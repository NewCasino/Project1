﻿Yapıkredi
