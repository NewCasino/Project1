Uttag av pengar direkt till ditt eKonto-konto