﻿Jackpottar