﻿Vänligen välj ett kort
