﻿/game/gamerules.jsp?game=viking&lang=sv