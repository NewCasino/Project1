Uttag direkt till ditt moneybookers konto