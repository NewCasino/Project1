Se alla alternativ!