﻿INSTADEBIT