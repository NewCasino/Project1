Uttag av pengar direkt till ditt AstroPayCard-konto