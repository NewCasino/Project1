﻿/game/gamerules.jsp?game=lrblackjackonedk&lang=sv