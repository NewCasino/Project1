Regler för Sportsbook