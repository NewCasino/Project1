<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktar  [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /> <br /> Din personliga insättning gräns är satt till $NEWLIMITAMOUNT$ $NEWLIMITPERIOD$. <br /> <br /> Du kan minska din insättningsgräns omedelbart i menyn Responsible Gaming på webbplatsen. <br /> <br /> Men om du vill öka din gräns, kommer det att ta 7 dagar innan den nya gränsen är aktiverad. 7-dagars perioden är till för att tillåta dig ompröva gränsen och byta vid behov. <br /> <br /> Tveka inte att kontakta oss om ni har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Kind Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kund Support Teamer </p>