Uttag direkt till ditt MasterCard kort.