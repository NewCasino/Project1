Öppnar kl.