﻿/game/gamerules.jsp?game=demolitionsquad&lang=sv