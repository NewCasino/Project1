﻿Väntande uttag
