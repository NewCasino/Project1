Debitera från {0} konto