Du har uppdaterat lösenordet