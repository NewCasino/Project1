﻿/game/gamerules.jsp?game=secretcode&lang=sv