﻿Bonus ej tillåten!
