Du får snart ett e-postmeddelande med ditt registrerade användarnamn.