﻿/game/gamerules.jsp?game=geisha&lang=sv