﻿<p>Kära kund,</p>
<p></p>
<p>Du måste acceptera  <a href="[Metadata:value(/Metadata/Settings.Terms_Conditions_Url)]" >Regler &amp; Vilkor </a> innan du kan spela.
</p>
<p>
 Tveka inte att kontakta våran kundstjänst om du har några frågor.
 </p>
 <p>
 <br />
 Tack så mycket, <br />
Kundtjänst
</p>

