Uttag från