﻿Trustly