﻿/game/gamerules.jsp?game=soccerslammini&lang=sv