﻿Ta ut pengar direkt till ditt bankkonto
