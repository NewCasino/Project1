﻿Välj Kreditkonto


