﻿Kings eller Bättre Serier

