﻿Klicka för att välja din bonus
