Glömt Lösenord