Länken är ogiltig eller har gått ut.