﻿Amerikansk Roulette
