﻿<!—Infoga loggan här -->
