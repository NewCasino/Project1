Fel, det här spelet kan inte spelas i helskärmsläge innan du har loggat in!