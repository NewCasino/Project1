Vänligen välj TLNakit konto