Andra banker