Laddning av saldon misslyckades.