jul