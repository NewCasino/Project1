﻿Skriv ut
