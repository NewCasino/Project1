﻿Kategory:
