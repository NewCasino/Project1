﻿Anmälningsavgift
