﻿Mina inställningar
