Ange förlustgräns