Oklart? klicka för att byta