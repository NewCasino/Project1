﻿Självexkludera i 1 år
