﻿Casino Poäng
