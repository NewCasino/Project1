Du har bytt lösenord