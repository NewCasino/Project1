Ett konto med samma detaljer är redan registrerat.