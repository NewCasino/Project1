Vänligen fyll i TC nummer