Användarnamn