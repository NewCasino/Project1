﻿Steg 2 / 2. 1 minut kvar...
