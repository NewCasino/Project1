﻿Gör ett uttag direkt från ditt UIPAS konto.
