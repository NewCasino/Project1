﻿Laddar...
