﻿Cancellation declined, subsequent tx issue.