Ta bort från Favoriter