penningbelöningar i hög takt