Skickat kl.