Kontoinnehavarens filial