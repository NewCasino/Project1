Israel shekel