Vänligen ange landet där du bor