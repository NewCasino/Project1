Gamla lösenordet