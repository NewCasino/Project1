(minus avgift)