Din anslutning har kopplats från eftersom du har uppnått tidsgränsen för din session.