Ange ditt lösenord!