﻿Du har ett väntande uttagsförfrågan. Vänligen vänta tills den bekräftas av vårt team. För mer information, vänligen kontakta vår livesupport.
