﻿WebMoney (från Moneta)