Transaktions-ID (valfri)