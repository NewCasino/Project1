Max. tillåten sessionstid (i minuter)