Rutnätsvy