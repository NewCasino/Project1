﻿Inbetalning med<span>{0}</span>
