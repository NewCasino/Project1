Moneybooker e-post