Aktiviteten har slutförts!