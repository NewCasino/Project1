Registrera dig