Hur fungerar det?