﻿Topp