Kompisens e-post