Du kommer inte kunna logga in på ditt vadslagningskonto under en period om 30 dagar för avkylning