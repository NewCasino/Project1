Din ändring av lösenordet lyckades.