Öppettider: