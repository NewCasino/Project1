﻿<p><span><strong>Villkor:</strong></span><br /><br />1. Det här erbjudandet gäller endast för ny registreade kunder hos Jetbull genom http://online.casinocity.com, den som gör sin första insättning på deras Jetbull Sportsbook konsto från och med den 1:a November 2012 till den 30:e November 2012.</p>
<p><br />2. Jetbull.com kommer att matcha första insättningen direkt gjord till Jetbull Sportsbook med en total bonus på 100% upp till maximalt &euro;50(eller motsvarande valuta)/$50/&pound;50. Both the deposit amount and bonus amount will be moved to bonus balance.</p>
<p>&nbsp;</p>
<p>3. Minumum insättningen första gången för första insättningsbonusen är på &euro;10(eller motsvarande valuta)/$10/&pound;10.</p>
<p>&nbsp;</p>
<p>4.För att kunna göra ett uttag av sin bonus, måst spelaren göra en total insats på deras insättning och insättningsbonus åtta (8) gånger med ett maximalbelopp &euro;50(eller motsvarande valuta)/$50/&pound;50, inom 15 dagar. Om satsingen är värd mer än &euro;50(eller&nbsp;motsvarande valuta)/$50/&pound;50, endast &euro;50(eller motsvarande valuta)/$50/&pound;50 kommer att räknas mot omsättningskravet.</p>
<p><br />5. Spelare kan kontrollera sin kvarstående omsättningskrav(en)(s) genomm att gå till&nbsp;<em>Mitt Konto -&gt; Aktivera Bonus</em>.</p>
<p><br />6. Om omsättningskravet inte är uppfyllt inom 15 dagar, kommer bonusar och vinster att bli förflyttade från kontot.&nbsp;</p>
<p><br />7. Dubbla satsningar eller plasterade satsningar på samma händelse kommer inte räknas mot satsningskraven.</p>
<p><br />8. Enkla, flera eller systemsatsningsbiljetter, både live och före live, med totala odds på 2.0 eller bättre är berättigade. För systemsatsningsbiljetter är minimum oddset på 2.0 gäller för selektion. Alla satsningar med läger odds än 2.0 kommer inte att räknas &nbsp;gentemo insatsen.</p>
<p><br />9. Detta erbjudande gäller för följande spelmarknader: Outright (Winner), Hästkapplöpning.</p>
<p><br />10. Våra bonusar är endast för våra hoppyspelare och Jetbull kan på samvete begränsa antalet kunder som får delta erbjudndet.</p>
<p><br />11. En bonus per kund, hushåll eller dator med delad IP är tillåtet.</p>
<p><br />12. Jetbull.com har rätten att beslag ta alla bonusar och/eller eventuella vinster om dåligt beteende uppvisas.</p>
<p><br />13. Jetbull.com  har rätten att stänga av spelare från det här erbjudandet om det finns anledningar att misstänka att erbjudandet missbrukas.</p>
<p><br />14. Detta erbjudande gäller inte för kunder från Belgien, Frankrike, Montenegro, Polen, Portugal, Ryssland, Serbien, Storbritanien, USA och Ukraina.</p>
<p><br />15. Spelare kan bli om bedda attvisa indetificaions dokument(KYC) för att bekräfta sin identitet. Vid felaktighet vid uppvisning av dokumenten kan det leda till att bonusar och/eller eventuella vinster tas bort.</p>
<p><br />16. Jetbull.com har rätten att stänga av denna bonus eller ändra villkoren när som helst.</p>
<p><br />17. Förutom ovannämda villkor, gäller det här erbjudandet under allmäna villkor.</p>
<p><br />18. Om händelse av en tvist uppstår ligger det slutliga beslutet hos Jetbull.com alltid.</p>
