<p>Hej $FIRSTNAME$,</p><p>Din insättning har genomförts.</p><p><span style="font-size: medium;"><strong style="color: #ff3366;">Vänligen klicka på "Refresh" knappen (inte web browserns refresh knapp) på sidan för att ladda sidan på nytt och se din balans.</strong></span></p><p>Om du har några frågor så tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>