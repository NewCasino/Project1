﻿Laddar...


