﻿Meddelande Sänt
