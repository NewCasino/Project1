<p>Hej $FIRSTNAME$,</p>Din insättning har nekats, vänligen kolla upp bankinformationen och försök igen senare.<p>Om du har några frågor gällande ditt kvitto var vänlig tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>