﻿Ogiltigt Konto ID.
