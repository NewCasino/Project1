Om det inte är fallet och du kom hit av en länk vi skickat till dig, länken kan vara utdaterad