Summa insatt till ditt {0} konto