﻿Let It Ride Serier
