﻿Självexkludera permanent
