﻿3-5 dagar