﻿Din väns fullständiga namn


