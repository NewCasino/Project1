[Metadata:value(/Metadata/Settings.Operator_DisplayName)], Ansvartfullt spelande