Ange mottagarens mobilnummer.