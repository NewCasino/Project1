Sätt in pengar