﻿Vänligen se bekräftelsekvitto på transaktionen
