﻿Underkänd anledning
