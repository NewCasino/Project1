Ta bort