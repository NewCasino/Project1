Visa spel i popularitetsordning