Sortera alfabetiskt