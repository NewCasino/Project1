Uttag av pengar direkt till ditt skrill-konto