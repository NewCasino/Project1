﻿eller
