Turkiet Banköverföring