Spelregler