﻿Hitta mer information om vårt belöningssystem
