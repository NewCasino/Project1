﻿Förnamn
