﻿Citizen ID
