﻿<ol>
 <li> <strong>Jag har glömt mitt användarnamn och lösenord, vad gör jag?</strong>
 <p>
Ett felaktigt angivet lösenord leder ofta till koden "kunde inte validera lösenord". Lösenord är skiftlägeskänsliga, kontrollera därför att du stängt av Caps Lock. Om problemet kvarstår, välj "glömt lösenord" så skickas ett nytt lösenord till den e-postadress som finns registrerat på ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto.
 </p>
 </li>

 <li> <strong>Vem ska jag kontakta om jag har frågor om mitt konto?</strong>
 <p>
Kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst
 <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">
 [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]
 </a>
 </p>
 </li>

 <li>
 <strong>Vad gör jag om jag inte vill använda mitt konto mer?</strong>
 <p>
För att stänga ditt konto [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst på
 <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">
 [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]
 </a>
 </p>
 </li>

 <li>
 <strong>Hur ändrar jag mitt lösenord?</strong>
 <p>
Du kan ändra ditt lösenord genom att använda "Glömt lösenord"
 <a href="/ForgotPassword" target="_blank">link</a>
 överst på alla [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] sidor.
 </p>
 </li>

 <li>
 <strong>Hur ändrar jag min registrerade e-postadress?</strong>
 <p>
För närvarande kan du inte ändra din e-postadress själv, men om du har goda skäl för ändring av e-postadressen, kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst för en ändring av dina kontouppgifter. Kontakta
 <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">
 [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]
 </a>
 </p>
 </li>

 <li>
 <strong>Hur kan jag kontrollera aktiviteten på mitt konto?</strong>
 <p>
Du kan kontrollera dina kontoaktiviteter genom att gå in på "Mitt konto" när du har loggat in,&nbsp; eller kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst för ytterligare information.
 </p>
 </li>

 <li>
 <strong>Kan jag ändra mitt användarnamn?</strong>
 <p>
Du kan inte ändra ditt spelarnamn när du har anslutit det till ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto. Detta för säkerhets skull eftersom ändring av spelarnamn kan störa systemets data och orsaka säkerhetslarm.
 </p>
 </li>

 <li>
 <strong>Vem kan jag kontakta om jag misstänker att jag har problem med mitt spelande?</strong> 
 <p>
Det är spännande, roligt och potentiellt vinstgivande att delta i onlinespel, för dem som väljer att spela. Men, [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] är medvetna om riskerna för spelmissbruk och följderna som det kan leda till för individen. Därför, [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] vidtar alla säkerhetsåtgärder för att säkerställa att våra produkter och tjänster endast används av personer som har laglig rätt att göra det. Spelare får under inga omständigheter spela om riktiga pengar om de inte uppfyller kraven om minimiålder på 18 år eller har uppnått lagenlig ålder för onlinespel i landet där de är stadigvarande bosatta.
 </p>
 </li>

 <li>
 <strong>Vad händer när min period har löpt ut?</strong>
 <p>
När tidsgränsen för din självuteslutningsperiod har löpt ut kan du kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst för att öppna ditt konto.
 </p>
 </li>

 <li>
 <strong>Hur kan jag utesluta mig själv?</strong>
 <p>
Du kan utesluta dig själv genom att gå in på ditt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] konto där du hittar fliken för självuteslutning och när du klickar på knappen Blockera mitt konto blir du automatiskt utloggad från [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] webbsidan. Därefter kan du endast logga in efter det att uteslutningsperioden som du valde har löpt ut.&nbsp; &nbsp;
 </p>
 </li>

 <li>
 <strong>Can I cancel it?</strong>
 <p>
 Du kan inte öppna ditt konto förrän tidsperioden som du valt för självuteslutningen har löpt ut.
 </p>
 </li>

 <li>
 <strong>Jag får inte svar på mina frågor när jag skickar e-postmeddelande till Kundtjänst?</strong> 
 <p>
Vi försöker besvara alla e-postmeddelanden till kundtjänst inom 24 timmar. Eftersom en del frågeställningar kräver mer detaljer och undersökningar kan svarstiden ibland variera beroende på frågans natur. Du får en bekräftelse via e-post från [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] när vi har tagit emot din fråga, för att meddela att vi arbetar på ett svar. Om du inte får en bekräftelse via e-post direkt efter det att du skickat din fråga, rekommenderar vi att du kontrollerar din Skräppost-korg. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] deltar inte i utskick av oönskade e-postmeddelanden men vissa aggressiva e-postfilter kan av misstag identifiera våra e-postmeddelanden som spam och behandla dem som sådana.
 </p>
 </li>
</ol>

<p style="text-align:right">
 <button type="button" onclick="window.print(); return false" class="button">
 <span class="button_Right">
 <span class="button_Left">
 <span class="button_Center">
 <span>Skriv ut</span>
 </span>
 </span>
 </span>
 </button>
</p>