﻿<!—Infoga logga här -->

