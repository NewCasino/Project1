﻿Fundsend