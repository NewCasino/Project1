﻿Vänligen skriv in mottagarens namn
