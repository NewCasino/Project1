Du har varit inaktiv för länge och din sittningstid har tagit slut. Av säkerhetskäl har du automatiskt blivit utloggad. Var vänligen tryck OK för att logga in igen.