﻿Säkerhetssvar
