Du kan inte spela förrän du klickat på länken i aktiveringsmailet. 