﻿Se gårdagens toppengaspelare
