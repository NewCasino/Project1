Uttag