Du har nu överfört pengarna.