﻿Ditt användar-ID måste bestå av minst 7 tecken
