﻿Video Poker
