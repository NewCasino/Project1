Användarnamnet måste innehålla mellan 4 och 20 tecken