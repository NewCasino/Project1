Uttag direkt till ditt CUENTADIGITAL konto