﻿You must sign in to your NETELLER account and accept the Terms and Conditions.