Spela nu