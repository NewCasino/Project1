Endast kvinnor