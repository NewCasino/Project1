Ange BOCASH-kod.