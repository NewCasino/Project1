E-postadress