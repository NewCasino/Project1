﻿Verifieringskoden har nu skickats till ditt mobilnummer. Kolla meddelandet.
