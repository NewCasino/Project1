﻿Registera Kort
