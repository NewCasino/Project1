Stäng helskärm