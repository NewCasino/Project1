﻿Popup
