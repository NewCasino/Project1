Växla vyn