Direkt banköverföring