Ange användarnamn och lösenord.