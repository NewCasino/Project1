﻿mgs-live-multispelare-roulette
