﻿Registrera ett Moneybookers-konto
