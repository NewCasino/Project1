﻿Insättning