Dölj fulla bord