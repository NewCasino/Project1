Ny e-postadress