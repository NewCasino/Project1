﻿IBAN är fel. Du får inte använda det angivna IBAN-numret.
