﻿Casino-plånbok FPP