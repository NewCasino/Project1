﻿Email är redan registrerad