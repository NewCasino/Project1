﻿ditt gamla lösenord här
