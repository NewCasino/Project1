﻿Beskrivning