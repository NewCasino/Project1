Uttag av pengar