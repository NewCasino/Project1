﻿Fyll i bankkod