Månad