Direktdebitering från ditt bankkonto