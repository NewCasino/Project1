﻿Enet Pokerbonus
