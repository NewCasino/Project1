﻿Ansvarsfullt spel
