﻿Din väns användarnamn


