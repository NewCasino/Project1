﻿Om oss
