Registreingen är klar