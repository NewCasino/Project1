Gör ett uttag direkt till ditt TrustPay konto