Slutsaldo