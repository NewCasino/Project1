[metadata:value(/Profile/_Index_aspx.Title)]