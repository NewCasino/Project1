﻿Överföring från ditt {0} konto