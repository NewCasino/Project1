﻿Självexkludering under 1 år
