﻿/game/gamerules.jsp?game=blackjackpntn&lang=sv