﻿Välj en checkbox!
