﻿Lösenordet måste innehålla minst 8 tecken