﻿/game/gamerules.jsp?game=subtopia&lang=sv