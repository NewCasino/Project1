﻿<p>Hej $FIRSTNAME$,</p>
<br />
<p>Användarnamn: $USERNAME$ </p>
<br />
Med detta mail vill vi bekräfta att din självexkluderingsperiod har nu avslutats. Du kan börja spela igen. 
<br />
<br />
Vänligen kontakta oss vid eventuella frågor på
<a href="mailto: [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]"> [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)] </a>
<p>&nbsp;</p>
<p>Med vänliga hälsningar,</p>
<p>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]  Kundtjänst </p>

