﻿3D animerat bordsspel 
