Beloppet passar inte för vald bonus