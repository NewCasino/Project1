Du kan snabbt göra en insättning från ditt Solo debet kort via Moneybookers till ditt spelkonto. Fyll i dina kortuppgifter via Moneybookers och när ditt kredikort kort är verifierat kommer din transaktion föras över till ditt spelkonto på en gång. 