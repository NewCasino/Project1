﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)], Ansvarsfullt spelande