﻿Sänder...


