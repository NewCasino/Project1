﻿Ditt UIPAS konto
