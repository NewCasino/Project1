﻿{0}d sedan