﻿vänligen ange koden
