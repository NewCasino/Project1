﻿Konto
