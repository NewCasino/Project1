﻿stäng detaljer
