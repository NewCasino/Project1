﻿This merchant does not support NETELLER (1-PAY) transactions.