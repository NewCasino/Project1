Avsändarens telefonnnummer