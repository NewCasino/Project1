Sydkorea Won