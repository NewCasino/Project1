﻿Filtrera specifika tillverkare...