Förnamn