﻿Favoriter