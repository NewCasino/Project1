Kontrollera att den valda valutan ovan är densamma som på din BOCASH-voucher.