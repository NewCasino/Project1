﻿Pay by SMS

