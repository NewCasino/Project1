Ange kortets utgivningsnummer.