﻿/game/gamerules.jsp?game=acescratch&lang=sv