TLNakit konto(n)