﻿System error