﻿[Metadata:value(.NegativeLimit_Style)]
<div class="NegativeLimitPanel">
<div class="NegativeLimitPopup">
    <div class="NegativeLimit_Content">
        <div class="NegativeLimit_Message_Text">
        </div>
    </div>
<a title="Close this popup now!" href="#" class="Close" onclick="$('.NactiveLimitPanel').hide();"> x </a>
</div>
</div>

