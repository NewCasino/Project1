﻿i-BANQ användar-MID lösenord är fel
