﻿Georgian Card - Leverantör av korthanteringstjänster.