Email är redan registrerad