Skapa ett lösenord