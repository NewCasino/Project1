Glömt lösenordet?