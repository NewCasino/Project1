﻿Säkerhets-ID/Autentiseringskod