﻿videokolikkopelit

