Du måste logga in för att se din tillgängliga bonus.