﻿Belopp som skall överföras till{0}
