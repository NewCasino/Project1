﻿SMS-kod