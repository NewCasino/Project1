Det upprepade lösenordet saknas