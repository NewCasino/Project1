﻿Lämna in
