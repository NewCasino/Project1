﻿Sport Matches
