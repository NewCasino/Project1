﻿Live Casino-bonus