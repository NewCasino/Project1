Spelinformation till {0}