﻿Förfallodatum : {0}