﻿/game/gamerules.jsp?game=allamerican5&lang=sv