﻿Jag vill inte sätta några gränser just nu
