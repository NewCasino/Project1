Bankens namn