﻿Din summan här
