﻿För många försök
