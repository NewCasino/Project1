﻿Gå Till: 
