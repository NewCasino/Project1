Referensnummer