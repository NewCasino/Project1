avgift taget