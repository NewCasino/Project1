Meddelanden