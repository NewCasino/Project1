﻿Trey Poker Serier
