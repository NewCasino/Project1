﻿/game/gamerules.jsp?game=frankenstein&lang=sv