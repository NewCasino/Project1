﻿Tillgängliga bonusar
