﻿Neteller(Ungern)
