Du kan inte spela det här spelet, komplettera din profil först.