Linjär vy