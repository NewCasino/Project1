﻿Ta ut direkt till din bank med Intelligent Payments
