Nästa