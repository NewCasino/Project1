Stad