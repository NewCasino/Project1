Registrera bankkonto