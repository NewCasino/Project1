Ta bort Favorit