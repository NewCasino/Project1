﻿Ukash Växel

