Gränsen har ändrats men den gäller fortfarande fram till utgångsdatumet. Nya beloppsgränser: