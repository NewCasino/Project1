Du kan inte göra en överföring till dig själv.