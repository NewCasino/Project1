﻿/game/gamerules.jsp?game=goldrushflash&lang=sv