Uttag av pengar direkt till ditt CASHU-konto