﻿Anmälningsavgit
