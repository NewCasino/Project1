Observera att du måste ha gjort minst en insättning för att kunna ta ut pengar från ditt konto.