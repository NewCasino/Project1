﻿Vänligen ange betalarens adress
