﻿Jag har en bonuskod
