nya spel