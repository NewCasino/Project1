Välj ett kort.