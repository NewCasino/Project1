﻿Notera: 

