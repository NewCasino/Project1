﻿Roulette Special