Växla mellan ikoner och lista.