﻿<P>Hej $FIRSTNAME$,</P>
<P>Välkommen till [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], vi vet att du kommer att trivas med att ta del av det roliga!</P>
<P>Ditt användarnamn är $USERNAME$, vänligen förvara detta på en säkert ställe så du håller en säker tillgång till ditt konto.</P>
<P>Om du inte redan har gjort det, så är det perfekt att ta del av våra välkomstförmåner. Du kan hitta alla erbjudande i vår kampanj sektion.</P>
<P> Om du har några problem med att signera upp dig, eller har några frågor till hos, tveka inte att höra av dig via <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>. Vi är här för att hjälpa och uppskattar din feedbback.</P>
<P>Med Vänliga Hälsningar ,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundservice</P>
