Elektronisk överföring