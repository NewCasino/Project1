Storbritanien , Pounds