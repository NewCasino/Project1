Välj landsnummer (prefix)