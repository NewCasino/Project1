﻿Jacks eller Better Video Poker Serier
