Uttag av pengar direkt till ditt CUENTADIGITAL-konto