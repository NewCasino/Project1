Ange ett positivt nummer.