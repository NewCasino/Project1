Gör en överföring enligt uppgifterna nedan.