﻿Trappa ned
