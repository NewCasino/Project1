﻿Voucher nummer måste vara 16 tecken.