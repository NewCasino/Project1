Kontrollsiffror