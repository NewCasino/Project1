﻿Ja, skicka mig mail med erbjudanden och viktiga nyheter. Jag vill också få SMS med exklusiva erbjudanden.
