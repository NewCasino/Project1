﻿Välkommen till
