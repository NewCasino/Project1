Betala med SMS