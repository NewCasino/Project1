﻿
<ol>
        
<li> <strong> Hur kan jag identifiera betalningar eller uttag till [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] ? på min bank/kreditkort uttalande </strong >
<p>
Alla insättningar och uttag som visas på antingen ditt kreditkort eller kontoutdrag kommer alltid åtföljas av en deskriptor som [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] kommer att nämnas . Detta gör att du kan hålla koll på dina insättningar till och uttag från platsen . </P >
</li >

<li> <strong> Kan jag använda mer än en betalnings metod ? </strong >
<p>
Ja du kan , men vi kan behöva underlag för eventuella förändringar i finansiella metoder . </P >
</li >

<li> <strong> Accepterar du kort från mitt land ? </strong >
<p>
Vi accepterar kort från alla lands utom USA , Turkiet och Frankrike . </P >
</li >



<li> <strong> Varför kommer inte din webbplats ta mitt kort ? </strong >
<p> Vissa kreditkort emittenter upprätthålla en regel som inte tillåter dig att göra direkta insättningar till spelsajter . Du kanske vill kontakta ditt kort för att diskutera denna fråga , eller prova någon av de e - wallet deponerar alternativ istället För ytterligare hjälp kontakta . [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] . Kundtjänst </p>
</li >


<li> <strong> Vad gör jag om mitt kort insättning får minskat eller förkastas ? </strong >
<p>
Ibland om du försöker sätta in en andra gång innan din senaste insättning har gått igenom , kan det räknas in i din 24-timmars och veckovis insättning gräns och därmed orsaka en insättning problem . Den vanligaste orsaken till detta att ske beror på felaktigt fylla i fälten i formuläret . Vänligen kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] kundservice för att få detta åtgärdat. Också Vissa kreditkort emittenter upprätthålla en regel som inte tillåter dig att göra direkta insättningar till spelsajter . Du kanske vill kontakta ditt kort för att diskutera denna fråga , eller prova någon av de e - wallet deponerar alternativ istället . </P >
</li >

<li> <strong> Kan jag använda mitt kort för att sätta in i min väns konto ? </strong >
<p> Du kan inte göra detta eftersom det anses vara en tredje part transaktion och under inga omständigheter tillåtet . </p >
</li >


<li> <strong> Jag har deponerats från fel kort av misstag - är det något jag kan göra </strong >
<p> Vänligen kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] Kundtjänst på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank"> [ Metadata : htmlencode (/Metadata/Settings.Email_SupportAddress ) ] </a > </p >
</li >


<li> <strong> Kan jag överföra pengar mellan konton ? </strong >
<p> Du kan inte föra över pengar mellan egna konton , men du kan överföra mellan Casino, Sport och Poker i ditt personliga konto . </p >
</li >


<li> <strong> Vad är ett IBAN-kontonummer? </strong >
<p> IBAN står för International Bank Account Number . IBAN används i internationella banktransaktioner tråd och gör att uttag av dina vinster lättare . </p >
</li >


<li> <strong> Vad är en CVC2 kod ? </strong >
<p> CVC2 är en akronym för " Card Verification Code " . Denna kod krävs som en säkerhetsåtgärd när man gör internationella telefonsamtal köp och betalningar internet med kreditkort . Denna kod består av tre siffror och återfinns på baksidan av ditt kreditkort .
</p >
</li >

</ol >

<p style="text-align:right">
    <button type="button" onclick="window.print(); avkastning false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span> Print </span >
                </span >
            </span >
        </span >
    </knappen >
</p >

























































 


 
 

 

 


 
 

 

 






Google Translate for Business:Translator ToolkitWebsite TranslatorGlobal Market Finder









Turn off instant translationAbout Google TranslateMobilePrivacyHelpSend feedback

