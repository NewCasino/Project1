﻿ditt bank konto
