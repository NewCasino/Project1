﻿Klassiset kolikkopelit
