﻿Din email här
