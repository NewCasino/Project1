Misslyckades