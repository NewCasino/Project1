﻿Taiwan