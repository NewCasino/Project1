Minsta poäng att göra anspråk på: