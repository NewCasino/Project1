﻿/game/gamerules.jsp?game=jackpot6k&lang=sv