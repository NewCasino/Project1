Peru Nuevo Sol