Populäritet