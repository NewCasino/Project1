Ungern forint