Du har för närvarande inga väntande uttag.  <br /><br />När du har ett väntande uttag här, har du möjlighet att cancelera transaktionen varvid dina medel omedelbart återvänder till ditt spelkonto. 