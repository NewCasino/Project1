﻿Jättipottipelit
