Populära