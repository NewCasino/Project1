﻿/game/gamerules.jsp?game=reddog&lang=sv