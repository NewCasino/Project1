﻿Få mail om nyheter och erbjudanden.
