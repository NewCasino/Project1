﻿Neteller(Australien)
