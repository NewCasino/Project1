﻿ditt nya lösenord här
