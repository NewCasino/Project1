Uttag direkt till ditt Switch/Solo kort.