﻿Demolition Squad™ är ett 5 reel, 4 rad och 40 bet line actionpakat högtenergi videoslot. Beskrivningen av demolition teams hårda arbetesdag på arbetet,  sloten erbjuder en stil i cartoongrafik med non-stop crew’s hard day at work, the slot offers cartoon style graphics with non-stop livlighet.

Demolition Squad™tar spelade spel till en exploderande levlar i Demolition Wild. Medan teamet arbetar på reels, spelare är förväntansfulla på att se det när två Wilds dyker upp på reels 2 och 4, alla symboler dyker upp mellan de två transformerade i Demolition Wild - ger chansen till en grundande vinst!

Players som förintar vägen till Free Spins upplever att Demolition Wilds fortsätter att ändra symbolder i wild. Men det som är mest spännanden är, vinster med Demolition Wilds med Free Spins är multiplicerade upp till x3.
