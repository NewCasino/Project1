Uppdatera din profil