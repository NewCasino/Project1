Uttag direkt till ditt PAGOFACIL konto