﻿Emailadressen finns redan i systemet
