<p>$USERNAME$,<br /><br />Tack för att du registrerat dig på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br />För din egen säkerhet vill vi påminna dig att verifiera din epost för att försäkra dig om att ditt konto fortsätter vara aktivt så att du kan fortsätta ta del av alla våra erbjudanden på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)].<br /><br /> Vänligen klicka på länken nedanför. Om det inte skulle fungera försök att kopiera länken och klistra in det i ett nytt fönster,<br /><br /><a href="$ACTIVELINK$">$ACTIVELINK$</a></p><br />Om du inte har registrerat dig hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], vänligen bortse från detta mail eller informera vår support  <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br /><p><br />Vänliga Hälsningar,<br />[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundservice teamet<br />