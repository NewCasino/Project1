Vänligen fyll i Ukash värde