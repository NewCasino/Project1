﻿Sportsbook
