Pengar överförs direkt till dit EcoCard kort