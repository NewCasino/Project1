Växla visning av spel från {0}