﻿/game/gamerules.jsp?game=cashbomb&lang=sv