Från mitt konto