﻿Verifieringskod

