﻿Ingen överföring har registrerats under den agivna tidsperioden.

