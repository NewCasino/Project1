Uttag direkt till ditt InstantDebit konto