Bonusar