Registrera kreditkort