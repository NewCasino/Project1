Uttag av pengar direkt till ditt InstantDebit-konto