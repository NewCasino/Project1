﻿/game/gamerules.jsp?game=casinoholdem&lang=sv