﻿Poker debet