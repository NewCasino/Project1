﻿Starta spel
