﻿Utfärda en IPS förbetald kupong och överför pengar till den nya kupongen.
