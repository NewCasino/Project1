Kompisens fullständiga namn