﻿/game/gamerules.jsp?game=fishyfortune&lang=sv