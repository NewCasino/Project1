Vi beklagar att inget av våra livebord är tillgängliga för dig. ({0}/{1}/{2})