﻿Venezuela