﻿Neteller(Schweiz)
