Välj period