Bonuskod