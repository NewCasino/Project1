﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Ditt uttag- IPS Token
