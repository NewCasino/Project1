Mottagarens namn