Spela LIVE Poker nu!