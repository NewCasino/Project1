Gäller fr.o.m.