Ogiltigt lösenord