Gränserna har ändrats, men fortfarande giltig fram till slutdatumet. Nya gränserna: