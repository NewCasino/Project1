Ogiltigt IBAN, du kan inte använda vårt exempel-IBAN.