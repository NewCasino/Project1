En 3 månaders självutslutningsperid