﻿Transaktion till spelare {0}