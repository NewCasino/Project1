Börsen måste börja med R / Z / E, följt av 12 siffror.