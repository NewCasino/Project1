﻿Lyckades