﻿/game/gamerules.jsp?game=retro-groovy60&lang=sv