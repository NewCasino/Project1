Konfiskera alla medel på förfallodagen