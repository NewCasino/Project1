﻿Tillgängliga Kort
