﻿Yandex (från Moneta)