﻿Klicka för att ange din bonuskod
