﻿Självexkludering permanent
