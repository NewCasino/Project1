Du har varit inaktiv för länge och din session har avbrutits. Av säkerhetsskäl har du loggats ut automatiskt.
Klicka på ok för att logga in igen.