﻿Bonus kod