﻿/game/gamerules.jsp?game=roulette2french&lang=sv