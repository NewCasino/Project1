﻿Mottagarens namn

