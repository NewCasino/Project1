Uttag av pengar direkt till ditt ePay-konto