﻿Intelligent Payments kopplar säljare och köpare i olika länder och hjälper till att sänka transaktionskostnader. 
