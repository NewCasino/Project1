Din hämtning av poäng lyckades.