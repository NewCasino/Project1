﻿Your payment card has been blocked