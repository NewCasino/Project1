﻿/game/gamerules.jsp?game=flowers&lang=sv