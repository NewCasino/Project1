Du måste logga in för att ta ut pengar.