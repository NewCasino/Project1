Kreditkort