﻿Heard And Mc Donald Islands