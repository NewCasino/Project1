﻿Säkerhetsfråga
