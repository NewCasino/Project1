Tack, din förfrågan kommer att bearbetas så snart som möjligt. 