År