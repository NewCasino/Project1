﻿Fyll i IBAN.