<p>Hej $FIRSTNAME$,</p><p>Du har begärt att din [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] e-mailadress ska ändras.</p><p>Av säkerhetsskäl måste vi be dig bekräfta din nya e-mailadress. För att göra detta, klicka på länken nedanför:</p><p><a href="$ACTIVELINK$">$ACTIVELINK$</a></p><p>Om denna länk inte svarar, kopiera och klipp in länken direkt i din webbläsare.</p><p>Om du inte vill ändra din e-mailadress, vänligen bortse från detta e-mail eller informera oss på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p>Vänliga hälsningar, <br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>