﻿Lösenord är inte samma
