Bank of Georgia är en kollektiv fullservicebank med erfarna bankirer och engagerad personal som är beredda att göra sitt yttersta för dig.