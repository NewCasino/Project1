﻿/game/gamerules.jsp?game=blackjackflash&lang=sv