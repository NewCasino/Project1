﻿Balans
