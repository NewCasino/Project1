﻿Ditt Ukash kort
