﻿Vänligen se till att din valuta är samma som BoCash vouchers valuta.
