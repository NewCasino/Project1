﻿i-BANQ användar-MID lösenord
