Ange innehåll.