Omgående