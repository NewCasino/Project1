﻿Credit till {0} konto.
