Ja tack, skicka mig anpassade erbjudanden via sms.