﻿Logga in på ditt befintliga [Metadata:value(/Metadata/Settings.Operator_DisplayName)] konto nu!