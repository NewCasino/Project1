Ange ditt lösenord