<p>Hej $FIRSTNAME$,</p><p>Du har använt en del av ditt Ukash kupongvärde och nedan finns dina nya detaljer för Ukash.</p><ul><li><strong>Ukash Kupong Nummer</strong>:$VOUCHERNUMBER$</li><li><strong>Ukash Kupong Summa</strong>:$VOUCHERAMOUNT$</li><li><strong>Ukash Kupong förbrukningsdag </strong>:$VOUCHEREXPIRYDATE$</li></ul><p>Om du har några frågor om din voucher tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet</p>