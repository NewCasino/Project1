﻿/game/gamerules.jsp?game=hrcstud2&lang=sv