﻿FPP Skattesatser
