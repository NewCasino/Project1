E-postadressen har existerat. Vänligen använd ett existerande konto!