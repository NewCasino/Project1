Välj titel