﻿Adress uppgifter

