﻿<p>Bästa $FIRSTNAME$,</p>
<br />
<p>Kontonamn: $USERNAME$ </p>
<br />
Med det här e-postmeddelandet bekräftar vi att din uteslutningsperiod nu har börjat och pågår till och med $EXPIRY_DATETIME$.  Under den här perioden kan du inte logga in på ditt konto. Vi meddelar dig via e-post när din självuteslutningsperiod är över.
<br />
<br />
Om du har frågor, tveka inte att kontakta oss på 
<a href="mailto: [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]"> [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)] </a>
<p>&nbsp;</p>
<p>Vänliga hälsningar,</p>
<p>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]  Kundtjänstteamet</p> 