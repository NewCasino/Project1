﻿Lösenordet måste innehålla bokstäver och siffror.
