﻿/game/gamerules.jsp?game=alienrobots&lang=sv