Land där du är stadigvarande bosatt