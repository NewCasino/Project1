﻿Belopp att dras från ditt konto.
