﻿/game/gamerules.jsp?game=cstudflash&lang=sv