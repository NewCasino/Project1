Betalningsmottagare