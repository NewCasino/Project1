﻿ny
