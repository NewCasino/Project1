﻿Oddskupong
