﻿Du kommer att omdirigeras till {0} sida för att fullfölja betalningen
