Ansökan