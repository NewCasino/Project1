﻿Tyvärr är denna sida inte tillgänglig.
