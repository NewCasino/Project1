Du måste bekräfta att du godtar regler och villkoren