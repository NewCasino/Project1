Du ansluter från en mobilenhet, vill du växla till mobilversionen?