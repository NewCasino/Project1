﻿Jag vill begränsa mitt spelande
