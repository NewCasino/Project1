Vinnare gratisspel