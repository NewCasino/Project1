﻿Din väns E-post
