Skapa en kod för att göra uttag från Bank of Georgia-bankomater.