Via menyn nedan kan du ange en gräns för maximal vadslagning per dag, vecka eller månad. När en gräns har angetts, får du ett bekräftelsemeddelande via e-post. Du kan minska din gräns när som helst via den här menyn. Men, om du vill ta bort eller öka din gräns tillämpas en väntetid på 7 dagar. Väntetiden ger dig tid att tänka över din ändring. Observera att den här vadslagningsgränsen endast gäller för Casino-spel.