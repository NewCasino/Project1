﻿<p>Hi $FIRSTNAME$,</p>
<p>Ditt uttag har slutförts.</p>
<p>
  <span style="font-size: medium;">
    <strong style="color: #ff3366;">Vänligen kontrollera saldot på ditt bankkonto.</strong>
  </span>
</p>
<p>
 Om du har några frågor tveka inte att kontakta  <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.
</p>
<p>
  Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team
</p>

