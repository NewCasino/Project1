﻿Cool-off anledning
