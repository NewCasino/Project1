Uttag av pengar direkt till ditt kort.