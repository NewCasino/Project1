Procentsatser