Banköverföringar