﻿/game/gamerules.jsp?game=footballcupmini&lang=sv