Mexiko,Peso