﻿Sätt gräns på omsättningen
