﻿/game/gamerules.jsp?game=diamondhunt&lang=sv