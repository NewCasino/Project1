Välkommen {0}@{1}, <a>Logga ut</a>.