﻿Spela på skoj
