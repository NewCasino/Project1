Se alla vinnare nu!