﻿<h2>Ditt konto har skapats.</h2>

<p>
	Genom att skapa detta konto har du också accepterat <a href="/TermsConditions">Terms and Conditions</a>, och att du vill bli kontaktad med kampanjerbjudanden via email. Om du önskar, kan du ändra det genom att gå in på <a href="/AccountSettings">Användarinställningar</a>.
</p>
<p>
	Du bör göra en inbetalning nu, så att du kan börja spela i vårt Casino och i vår sportsbook!
</p>
