Transaktionshistorik