﻿andra-spel
