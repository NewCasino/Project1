Uttag direkt till ditt EPS konto