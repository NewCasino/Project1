Kampanjkoden har gått ut.