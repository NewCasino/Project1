﻿Kontakta Oss
