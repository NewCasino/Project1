﻿PayCard status was not changed