﻿<ol>

    <li> <strong>Vad är systemets minimikrav för att spela på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]?</strong> 
        <p>
            <ul>
                <li>
                    Windows - Intel Pentium processor (Pentium II eller högre rekommenderas) 64mb ram.
                </li>
                <li>
                    Macintosh - Power Macintosh Power PC processor (G3 eller högre rekommenderas) 64mb ram.
                </li>
                <li>
                    Viktig information till Apple Mac-användare - Nuvarande version av Casino kanske inte fungerar som avsett på ett Mac-system från Apple och stöds inte för närvarande.
                </li>
                <li>"FLASH" 10 eller högre</li>
                <li>
                    [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] är kompatibel med de flesta Windows operativsystem (Windows 2000, XP, Vista och 7).
                </li>
                <li>Internet Explorer-versioner lägre än 7 stöds inte.</li>
            </ul>
        </p>
    </li>

    <li> <strong>Vad händer om min anslutning bryts?</strong>
        <p>
            Alla spelomgångar lagras säkert i våra servrar och efter eventuella avbrott i anslutningen kan du enkelt logga in på ditt konto igen och se resultaten för alla händelser eller spelade spel. Detsamma gäller casinot, om en spelomgång inte hade slutförts ska den återupptas nästa gång du loggar in på spelet igen. Upplever du fortsatta problem, "klicka här" för att chatta med personalen på vår Kundtjänst.
        </p>
    </li>

    <li>
        <strong>Vilken programvaruleverantör använder ni?</strong>
        <p>
            Programvaran för vår sportbok är Oddsmatrix, Casinot har Net Entertainment och vår Poker använder Cake.
        </p>
    </li>

    <li>
        <strong>Varför kan jag inte ansluta till spelservern?</strong>
        <p>
            Kontrollera din internetanslutning och om problemet kvarstår, kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst.
        </p>
    </li>

    <li>
        <strong>Varför kan jag inte logga in på mitt konto?</strong>
        <p>
            Kontrollera att du använder rätt "lösenord" och "namn" på ditt konto, om problemet kvarstår kontakta [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst.
        </p>
    </li>

    <li>
        <strong>Webbsidan är mycket långsam, vad kan jag göra för att snabba upp den?</strong> 
        <p>
            Om du upplever att anslutningen är långsam, tänk på följande: Om du har flera webbläsare öppna, använder musikprogram eller laddar ned filer kan dessa göra datorn och/eller internetanslutningen långsammare. Det kan även lagga hos din lokala internetleverantör. Anslutningen kan även bli långsammare om du delar internetanslutning inom ditt hushåll och ditt lokala område.
        </p>
    </li>

    <li>
        <strong>Jag har inget ljud.</strong>
        <p>
            Kontrollera att du har ett giltigt ljudkort och att dina högtalare inte har stängts av. Kontrollera att du har ljudnivån inställd via [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] fliken "Alternativ". Chat-fliken nederst i högra hörnet på skärmen har en "Alternativ"-knapp där du kan välja "alla", "endast varningar" eller "tyst".
        </p>
    </li>

    <li>
        <strong>Har ni en MAC-version?</strong>
        <p>
            Tyvärr, vi kan för närvarande inte erbjuda någon version av programvaran som är särskilt framtagen för MAC. Många av våra användare har dock lyckats koppla in en PC-emulator för att kunna spela våra spel. Besök vår nedladdningssida för ytterligare information.
        </p>
    </li>

    <li>
        <strong>Varför är mitt spel så långsamt?</strong>
        <p>
            Kommunikationen mellan din maskin och våra servrar har optimerats för snabbast möjliga respons. Om du upplever att ditt spel är långsamt, kan det bero på två saker: 1. Spelarna vid bordet tar lång tid på sig att agera när det är deras tur. 2. Du kanske inte har en bra internetanslutning.
        </p>
    </li>

</ol>
<p style="text-align:right">
    <button type="button" onclick="window.print(); return false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span>Print</span>
                </span>
            </span>
        </span>
    </button>
</p>