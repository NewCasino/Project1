﻿PågåendeDebit