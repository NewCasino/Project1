Visa spel i en lista