﻿{0} tillgängliga
