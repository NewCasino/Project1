Din väns konto är blockerat