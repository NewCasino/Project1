﻿Cool-off för 3 månader
