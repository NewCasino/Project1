Vänligen välj mottagarens födelsedatum