﻿Hemsidans utseende och känsla
