﻿Välj kreditkort
