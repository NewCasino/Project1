Adressuppgifter