﻿Registrera