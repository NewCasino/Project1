﻿<h2> Ditt konto har skapats. </h2>

<p>
Genom att skapa detta konto har du också godkänt användarvillkoren <a href="/TermsConditions"> villkor </a>, och att du vill bli kontaktad för kampanjerbjudanden via e-post. Om du vill, kan du ändra det genom att gå <a href="/AccountSettings"> Användarinställningar </a>.
</p>
<p>
Du bör göra en insättning nu, så du kan börja spela på vårt casino och börja satsa på vår sportsbook!
</p>
