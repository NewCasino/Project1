﻿/game/gamerules.jsp?game=tribble&lang=sv