Skrill-konto