Ändra maxsumma