﻿OS spel
