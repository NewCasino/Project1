Uttag av pengar direkt till ditt UkashHosted-konto