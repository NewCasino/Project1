﻿Förnamn måste anges
