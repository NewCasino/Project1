﻿/game/gamerules.jsp?game=hrtxsholdem&lang=sv