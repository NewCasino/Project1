Laddar saldon...