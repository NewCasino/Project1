Ange ämne.