﻿Gör ett uttag direkt till bank via DengiOnline

