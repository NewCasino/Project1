Du kom troligast till denna sida av misstag.