﻿Voucherkod
