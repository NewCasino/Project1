﻿TXS Hold'em Serier
