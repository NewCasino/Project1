Registreingen