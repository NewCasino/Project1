﻿<p>Hi $FIRSTNAME$,</p>
Din insättning nekades, vänligen kontrollera bankinformationen och försök igen senare.
<p>Om du har några frågor angående ditt kvitto tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p>
<p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>



