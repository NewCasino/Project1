﻿Överföring
