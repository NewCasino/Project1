﻿Jacks eller Better I
