Välj din bank