Obegränsat antal säten