﻿Poker kredit