﻿<img src="//cdn.everymatrix.com/_casino/3/388A34DF99ECFA9F5B01EA8EE19B811B.jpg" />
