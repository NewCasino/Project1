﻿<ol>

    <li> <strong>Jag har laddat ner programvaran - var är den?</strong>
        <p>
            When the [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Poker software has been successfully installed to your computer, a [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Poker icon will appear on your desktop. Simply double-click on this icon to launch the poker software and you'll be taken immediately to our Game Lobby.
        </p>
    </li>

    <li> <strong>My password isn't being accepted?</strong>
        <p>
            Entering an incorrect password can often result in an 'unable to validate password' code. As passwords are case sensitive, check to ensure your Caps Lock is off. If your troubles persist, select the 'forgot password' button and a new password will be issued to the e-mail address as listed on your [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] account.
        </p>
    </li>

    <li>
        <strong>Can I change my nickname?</strong>
        <p>
            [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Poker allows players the ability to change their Player ID (name appearing at the poker tables) every 7 days. To do this, please visit the 'My Account' tab when logged on to the [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Poker software.
        </p>
    </li>

</ol>

<p style="text-align:right">
    <button type="button" onclick="window.print(); return false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span>Print</span>
                </span>
            </span>
        </span>
    </button>
</p>