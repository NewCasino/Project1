﻿Direkt banköverföring (med GPaySafe)
