Ange ett telefonnummer med 7 till 30 siffror