﻿/game/gamerules.jsp?game=megajoker&lang=sv