Ange kortets säkerhetskod.