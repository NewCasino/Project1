Ange Ukash-nummer