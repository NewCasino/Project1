Georgien Lari