﻿scratch-cards