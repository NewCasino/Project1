﻿/game/gamerules.jsp?game=lrhilo2-3c&lang=sv