﻿Betalarens adress
