Uttag av pengar direkt till ditt EUTELLER-konto