Har du inget NETELLER-konto? Klicka <a href="/Deposit/NetellerQuickRegister">här</a> för att registrera ett.