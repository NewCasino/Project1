﻿Jackpott
