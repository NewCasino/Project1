Din kompis konto är inaktiverat.