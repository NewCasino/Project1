﻿<p>Hej $FIRSTNAME$,</p>

<p>Det här är en bekräftelse på att din e-postadress på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] har ändrats enligt din begäran.</p>
<p>Om du inte har begärt ändring av din e-postadress, meddela omedelbart vår kundtjänst på 
<a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>
</p>

Vänliga hälsningar, 
[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänst