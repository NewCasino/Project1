Din anslutning har kopplats från eftersom din IP-adress har ändrats sedan din senaste inloggning.