Hjälp