Skattekod