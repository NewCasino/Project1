﻿Transaktions-ID