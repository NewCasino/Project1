﻿i-BANQ användar-MID
