﻿Pöytäpelit
