Du spelar i underhållningsläge. För att spela med riktiga pengar, logga in först.