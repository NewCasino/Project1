[Metadata:value(/Metadata/Settings.Operator_DisplayName)] – Din insättning har accepterats.