Det här fältet är obligatoriskt