Åtgärden lyckades!