Ja, skicka mig e-postmeddelanden om nyheter och erbjudanden.