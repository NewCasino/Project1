Uttag direkt till ditt PRZELEWY konto