﻿/game/gamerules.jsp?game=luckyeight&lang=sv