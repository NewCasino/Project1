﻿/game/gamerules.jsp?game=scratchticket&lang=sv