Fyll i användarnamn och lösenord