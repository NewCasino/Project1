﻿/game/gamerules.jsp?game=champion&lang=sv