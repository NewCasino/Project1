Vänligen se till att du noterat dina ändringar då du inte kan gå tillbaka till detta fönster. 