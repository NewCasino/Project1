﻿Referens ID
