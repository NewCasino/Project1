﻿Okt