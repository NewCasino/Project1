﻿Payment declined. Please activate your default Payment Method and try again.