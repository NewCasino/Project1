Mottagarens födelsedatum