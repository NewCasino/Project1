Vänligen fyll i ämne. 