ange din 1-Tap-gräns