Vänligen ange ditt svar på din säkerhetsfråga