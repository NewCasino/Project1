Utfärda ett kort