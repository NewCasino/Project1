Sortera spelen