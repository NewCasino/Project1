﻿/game/gamerules.jsp?game=luckyeightsafari&lang=sv