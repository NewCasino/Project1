OBS!