Betala per telefon (Portugal)