﻿Skriv in ditt användarnamn
