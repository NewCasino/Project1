Ange betalningsmottagare.