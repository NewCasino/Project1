﻿Voucher nummer är obligatorisk.