Du kommer få ett mail med instruktioner om hur du byter lsöenord