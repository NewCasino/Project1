﻿Överför till en vän

