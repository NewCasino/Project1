﻿Vänligen välj ett spelkonto.
