﻿Sammanslagna pokerturneringar
