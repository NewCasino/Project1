Ange SWIFT.