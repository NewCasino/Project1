﻿<p>Bästa $FIRSTNAME$,</p>
<br />
<p>Kontonamn: $USERNAME$ </p>
<br />
Med det här e-postmeddelandet bekräftar vi att din uteslutningsperiod är över och alla kontofunktioner är nu aktiverade.
<br />
<br />
Om du har frågor, tveka inte att kontakta oss på 
<a href="mailto: [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]"> [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)] </a>
<p>&nbsp;</p>
<p>Vänliga hälsningar,</p>
<p>[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Kundtjänstteamet</p>