Free HTML för innehållet är redigeringsbart i CMS Console.