﻿Kontoinformation
