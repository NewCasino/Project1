﻿Bank
