Gå till toppen