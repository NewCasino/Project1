﻿Bankkontonummer
