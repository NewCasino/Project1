﻿SNS Bank
