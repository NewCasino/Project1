Fler filter