﻿[metadata:value(/Metadata/Settings.Operator_DisplayNameShort)]
