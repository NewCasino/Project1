Inaktivera bakgrunden