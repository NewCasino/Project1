Daglig gräns (per dag)