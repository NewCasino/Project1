﻿Anledning till nedtrappning
