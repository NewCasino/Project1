Uttag av pengar direkt till ditt WebMoney-konto