﻿Välj valuta
