﻿Din födelsedata här (DD/MM/YYYY)
