Ange ditt ID-nummer.