﻿Wild Rockets
