﻿Neteller(Norge)
