Kortnummer behövs