﻿Adjustment declined - no reference ID