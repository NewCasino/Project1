﻿[metadata:value(/Metadata/Settings.Operator_DisplayName)] Mobile

