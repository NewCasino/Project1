Allmänna frågor om casino