﻿Pris pool 
