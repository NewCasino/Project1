Välj önskat öppningsläge för spelet här, inklusive inline / popup / ny sida och helskärm.