Öppnar spelet överlappande.