﻿/game/gamerules.jsp?game=lrroulettemini&lang=sv