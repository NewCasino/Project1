Platsernas status: