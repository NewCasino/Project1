<p>Hej $FIRSTNAME$,</p><p>Din insättning har lyckats.</p><p><span style="font-size: medium;"><strong style="color: #ff3366;">Vänligen tryck på “Uppdatera” knappen(INTE webbläsarens uppdateringsknapp) på sidans huvudfält för att uppdatera saldot.</strong></span></p><p>Om du har några frågor var vänligen tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Hälsninar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>