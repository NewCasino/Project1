﻿Poker saldo

