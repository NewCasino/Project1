Vänligen ange ditt mobilnummer