Du kan inte logga in eftersom du är från ett som omfattas av restriktioner.
Har du problem, kontakta kundtjänst.