Address rad 2