﻿Banköverföring till bankkonto i Turkiet kan endast skötas i EUR eller USD, vänligen se till att din bank accepterar banköverföringar I EUR eller USD
