﻿Mitt Konto

