Insättning