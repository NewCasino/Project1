Du är inte berättigad att göra en insättning.