﻿<p>Kära $FIRSTNAME$,</p>
<br />
<p>Kontonamn: $USERNAME$ </p>
<br />
Detta mail är en bekräftelse på att din självexkluderingsperiod has slutat och att ditt konto kommer aktiveras den $EXPIRY_DATETIME$.
<br />
<br />
Tveka inte att kontakta oss om du har några frågor eller funderingar på<a href="mailto: [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]"> [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)] </a>
<p>&nbsp;</p>
<p>Vänliga hälsningar,</p>
<p>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]  Kundtjänst</p> 

