Ange din e-postadress.