﻿Nätsluss
