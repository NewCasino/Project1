﻿Spel RTP
