﻿Din identitet måste verifieras innan du kan göra en överföring.
