Mitt favoritlag?