Landsnummer (prefix)