<p>Kära $USERNAME$,<br /></p><br />Syftet med detta e-mail är att bekräfta att ditt konto nu är install på självutslutning.<br /><br />Du kommer inte längre kunna logga in på ditt konto.<br /><br />Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><br /><br /><p>Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>