﻿Sidans design och upplevelse
