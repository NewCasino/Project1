Påminn mig inte igen