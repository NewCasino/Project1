Din address måste innehålla minst 2 tecken