﻿Tackar för din tid med oss!
