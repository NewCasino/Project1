﻿/game/gamerules.jsp?game=allamerican25&lang=sv