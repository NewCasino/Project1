Dagliga toppvinnare