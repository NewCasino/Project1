Visa spel i populäritetsordning