Spela {0} med riktiga pengar!