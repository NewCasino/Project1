﻿Thief™ är ett 5-reel, 25 bet video slot maskin Expanderar Wild symboler, regulära Gratis Spinns och Adrenalinfyllda Gratis Spinns med tillägg bar sympol; Diamant symbolen.
