Välj mottagarens födelsedatum.