﻿Kvitto
