﻿/game/gamerules.jsp?game=horserace&lang=sv