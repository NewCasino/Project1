Ange TC-numret.