Klicka <a href="http://www.playcoins.net/" target="_blank" title="Play Coins">här</a> för att köpa mynt. 