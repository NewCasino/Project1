Datum och tid