﻿OBS! Du kan endast byta in jämna <span class='messageHighlight'>{0}</span> poäng för 
<span class='messageHighlight'>{1} {2}</span>, resterande poäng sparas på ditt FPP-konto.