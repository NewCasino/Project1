﻿Intelligent Payments
