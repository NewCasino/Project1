﻿Debit från {0} konto.
