Skrill e-postadress