Bekräfta mobilnummer