﻿Euro600