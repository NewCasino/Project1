﻿<p>Kära $FIRSTNAME$,</p>
<br />
<p>Kontonamn: $USERNAME$ </p>
<br />Detta mail är en bekräftelse på att din nedträppningsperiod har slutat och alla funktioner har nu aktiverats på ditt konto.
<br />
<br />Tveka inte att höra av dig till oss om du har några frågor eller funderingart 
<a href="mailto: [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]"> [Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)] </a>
<p>&nbsp;</p>
<p>Vänliga hälsningar,</p>
<p>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]  Kundtjänst</p> 
