Lojalitet belönas på Guts Casino - och med belöning menar vi rena pengar! 