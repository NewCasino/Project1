﻿Tillbaka



