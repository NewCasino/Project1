﻿Batch status '{0}' can not be updated on '{1}'