Din kompis identitet är inte verifierad.