﻿Skickar

