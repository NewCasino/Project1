﻿/game/gamerules.jsp?game=relicraiders&lang=sv