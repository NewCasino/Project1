Avsändarens TC-nummer kan inte vara tomt.