﻿Att dras från {0}
