Ange ett belopp som ska överföras.