﻿Captcha är felaktigt, vänligen prova igen
