De kommande 30 dagarna