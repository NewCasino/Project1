﻿/game/gamerules.jsp?game=thrillspin&lang=sv