﻿Inloggningen ej tillåten!
