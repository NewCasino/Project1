Betala per telefon (Tyskland)