Din e-postadress