﻿Vänligen ange ett korrekt datum
