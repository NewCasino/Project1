﻿/game/gamerules.jsp?game=jackandbeanstalk&lang=sv