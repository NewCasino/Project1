Överför alla