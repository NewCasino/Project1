﻿Maxlängd för beskrivningen är 100 tecken
