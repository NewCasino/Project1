﻿/game/gamerules.jsp?game=fruits&lang=sv