Välj befintligt konto