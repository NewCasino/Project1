﻿Nummer
