Ukash värde