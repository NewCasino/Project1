﻿Sic Bo