Vadslagningskrav förlopp