Hem Bonus