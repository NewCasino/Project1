Välj konto