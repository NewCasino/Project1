Danmark, Kroner