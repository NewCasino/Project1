Ditt mobilnummer har redan registrerats.