Registrera ett TLNakit-konto