Variabler