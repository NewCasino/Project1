﻿Neteller(Nederländerna)
