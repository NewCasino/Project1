Snabbinsättning