Agentens kod