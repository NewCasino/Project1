Dotterbolag