﻿Du måste bekräfta att du är 18 år eller äldre och godkänna regler och villkor
