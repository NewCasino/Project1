﻿Inloggningen misslyckades. Du har valt att självexkludera dig från spel till {0}. Vänligen kontakta supporten då.

