﻿Hoppa over 
