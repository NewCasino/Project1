﻿Kasinobonus
