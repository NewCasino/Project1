﻿/game/gamerules.jsp?game=deadoralive&lang=sv