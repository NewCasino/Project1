﻿<ol>
        
<li> <strong> Vilka är de lägsta och högsta insats tillåtet ? </strong >
<p> Maxinsats varierar beroende på evenemanget . Om du försöker att placera satsningar som överstiger den maximala gränsen , kommer du att få ett meddelande som talar om det högsta belopp som du har rätt att satsa på det valet . Vi har inte en minsta insats begränsning . <p>
</li >

<li> <strong> Vad är singelspel och flera satsningar ? </strong >
<p> Singelspel innebär bara ett val , en multipel insats kräver mer än en . Ju fler val du länkar ihop i en multipel ( t.ex. alla hem lag i en omgång av Premier League ) , desto mer kan du vinna - men det är naturligtvis mycket svårare <p>
</li >

<li> <strong> Hur många val kan en flerfaldig satsning innehålla ? </strong >
<p> maximala antalet val vi gör i en multipel insats är 10 . <p>
</li >

<li> <strong> Hur handikapp vadslagning arbete ? </strong >
<p> För detaljerade förklaringar av handikapp vadslagning ( 1x2 med handikapp och asiatiska handikapp ) , besöka Betting Förklaring avsnittet här . <p>
</li >

<li> <strong> Vad händer om en match skjuts upp ? </strong >
<p> Kontrollera reglerna för denna sport . Vissa sporter kräver att matchen ska spelas på samma dag för att spelen ska gälla , kan satsningar inom andra sporter vara öppna tills matchen är klar eller officiellt övergivits . <p>
</li >

<li> <strong> Varför har mitt vinnande spel ännu inte betalats ? </strong >
<p> [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] kräva officiella resultat som skall deklareras innan marknaderna kan lösas . Ibland källor på nätet som live score platser kan vara felaktig så avveckling kan fördröjas tills resultaten kan bekräftas . <p>
</li >

<li> <strong> Jag har ändrat mig , kan jag avboka min insats ? </strong >
<p> Nej När du har bekräftat din insats och det har accepterats av vår server , kan spel inte annulleras . <p>
</li >

<li> <strong> Var kan jag hitta en förteckning över mina spel? </strong >
<p> din vadslagning och historier transaktionen kan hittas under " Mitt sportbetting konto " när du loggar in på [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] hemsida <p> .
</li >

<li> <strong> Varför är vinster beräknas på olika sätt på brittiska odds ? </strong >
<p> Vid beräkning vinster , använder vi decimal ( EU ) odds som de är mest korrekta . UK och US odds endast för visning ändamål som vissa decimalodds inte korrelerar till ett enkelt bråk . <p>
</li >

<li> <strong> Betting blir beroendeframkallande för mig , vad kan jag göra ? </strong >
<p> Betting med [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] bör vara ett roligt tidsfördriv för alla , men för en liten minoritet av människor , kan det bli beroendeframkallande och skapar problem . Information om spelberoende kan hittas via Ansvarsfullt spelande . <p>
</li >

</ol >
<p style="text-align:right">
    <button type="button" onclick="window.print(); avkastning false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span> Print </span >
                </span >
            </span >
        </span >
    </knappen >
</p >
