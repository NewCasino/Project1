﻿/game/gamerules.jsp?game=jacksorbetter25&lang=sv