﻿Information


