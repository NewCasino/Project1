﻿Logga in med
