﻿Neteller(Sydafrika)
