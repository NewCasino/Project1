Belopp som ska debiteras från {0} konto: {1} {2}