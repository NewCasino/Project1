﻿Självexkludering
