Ditt användarnamn innehåller otillåtna tecken