Välj ett användarnamn