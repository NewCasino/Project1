﻿Skicka
