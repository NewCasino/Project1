Sön