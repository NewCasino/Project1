Klicka här