Obegränsad