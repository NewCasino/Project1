Debeitera från {0} konto