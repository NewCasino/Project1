Ange IBAN.