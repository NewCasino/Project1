Ogiltigt kortnummer