Bonuskoden har aktiverats!