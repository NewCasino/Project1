Välj land