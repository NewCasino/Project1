﻿Bekräfta
