﻿TC-nummer