I linje