Lägg {0} till i Favoriter