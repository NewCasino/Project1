﻿Gör ett uttag från ett annat konto
