Välj ett Skrill-konto.