﻿Anledning till att du är otillfredställd
