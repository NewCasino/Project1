Ange ditt telefonnummer