Uttaget kommer att behandlas så snart som möjligt.