﻿Sätta in
