Bearbetar