﻿Du måste välja en av tillgängliga alternativ
