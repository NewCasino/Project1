﻿Maxlängden för fältet avsedd för efternamn är överskriden
