﻿Bordspel
