﻿Ge ut en Ukash förbetald kupong och överföra pengar till den nya verifikationen.
