Förfallodatum