Du har uppdaterat ditt lösenord