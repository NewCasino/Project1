﻿Alternativ för uttag
