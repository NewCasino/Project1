En 30 dagars självutslutningsperiod