Ta bort {0} från favoriter