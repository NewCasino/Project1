﻿Land Blokerat

