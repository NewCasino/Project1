﻿PayKwik (By MoneyMatrix)