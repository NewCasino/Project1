Ange vadslagningsgräns