﻿Klassiska Automater
