Gränser