﻿Populärt
