﻿Registrera Dig

