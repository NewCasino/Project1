﻿Spelutvecklingsbonus
