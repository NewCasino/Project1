﻿Notering: Du kan endast byta i omgångar <span class='messageHighlight'>{0}</span> poängen för 
<span class='messageHighlight'>{1} {2}</span>, de kvarstående poäng kommer att finnas kvar i ditt FPP konto.
