﻿Neteller(Estonien)
