﻿Jacks eller Better II
