﻿Pågående Utbetalning
