﻿/game/gamerules.jsp?game=thvideopokerjob&lang=sv