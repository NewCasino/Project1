Lör