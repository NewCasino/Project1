﻿Click2Pay