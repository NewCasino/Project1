﻿/game/gamerules.jsp?game=ghostpirates&lang=sv