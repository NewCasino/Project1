Uttag direkt till ditt CASHU konto