﻿Alla spel
