Välj