Tomt fällt: [ $FÄLT$ ]