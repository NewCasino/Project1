﻿Utfärda en IPS förbetald kupong och överföra pengar till den nya verifikationen.
