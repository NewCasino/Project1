Kompisöverföring