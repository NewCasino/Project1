Lö