﻿Beloppet är utanför gränserna


