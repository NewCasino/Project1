Säkerhet