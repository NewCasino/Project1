﻿Självexkludering under 5 år
