Ange tecken.