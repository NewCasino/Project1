﻿Namn
