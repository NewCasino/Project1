Till konto