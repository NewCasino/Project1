﻿Kontonummer