Typ av gräns