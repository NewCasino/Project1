De kommande 3 månaderna