﻿Från mitt konto


