Vadslagningsgräns