﻿poytapelit
