Emailet kunde inte skickas, försök igen.