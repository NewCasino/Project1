Jag bekräftar att jag är 18 år eller äldre och har redan accepterat era 