Nordea Solo Finland