Jag önskar ta emot alla tillämpliga bonusar.