﻿<p>Lojalitet har belöningar på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kasino - och genom belöningar menar vi hårda kontanter!
</p>
<br/>
<strong>Earning Casino Frequent Player Points</strong>
<p>
När du spelar kasinospel på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] med riktiga pengar,
du tjänar Kasino poäng på alla spel. Dessa poäng kan omvandlas till kontanter när du vill så länge du har ett saldo på minst 200 poäng eller mer. 
</p>
<br/>
<strong>View and Claim Points</strong>
<p>
Du kan
alltid övervaka dina Kasino Poäng-saldo på kasino sidan, och kom ihåg,vid [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] vi handlar om fair play, så tjänade poäng ska aldrig upphöra.. 
För att omvandla dina Ckasino poäng to money, till pengar, bara klicka på Lås knappen nedanför Kasino Poäng-saldon. Varje 100 poäng betalar € 1 och dessa medel är ska direkt till ditt konto.Om du har valt en annan valuta för ditt kasinokonto, du kommer att få motsvarande 1 € per 100 Poäng betalas i önskad valuta. 
</p>
<br/>
<strong>Earning Points </strong>
<p>Spel
genererar Kasino Poäng vid olika hastigheter.
 Se på regler och villkor nedan för att se hur många poäng du tjänar visst du spelar dina favoritspel.. 
Hastigheten är uttryckt i procent, vilket innebär hur mycket av ett casino poäng du tjänar varje gång du satsar € 1. Och naturligtvis, alla spel räknas, även om du satsar mindre än € ​​1. 
Till exempel, en av våra populära videoslots, Gonzo's Quest, tjäna i en takt på 20%. Detta innebär att om du satsar € 10, kommer du att tjäna 2 Kasino Poäng. 
</p>
<br/>
<strong>S</strong>
<p>
Speciella kampanjer</strong>
<p>Kolla efter våra unika Cash Rewards kampanjer. Ibland ökar vi skattesats för vissa spel under en tidsperiod. Kolla in nyheterna på kasino sidan, för spel som tjänar ännu högre takt. 
</p>
<br/>
<strong>Terms & Conditions</strong>

<ol class="fpp_termsconditions_list">
<li>Alla kunder tjänar Kasino Frequent Player Poäng visst man spelar kasinospel med riktiga pengar. </li>
<li>Minst 200 Kasino Poäng krävs för att omvandla poäng till pengar. Var 100 Kasino Poäng konverteras till € 1 (eller motsvarande valuta). Vid konvertering, förblir överblivna punkter som inte spenderas i kundens Kasino Poäng-saldon. </li>
<li>Spelets hastighet uttrycker hur många procent av insats Kasino Poäng genererar på € 1 (eller motsvarande valuta). </li>
<li>Alla spel i kategorierna Video Slots, Classic Slots, Progressive Slots, Scratch Cards och andra spel genererar poäng i en takt på 20%, alla Video Pokers och Bord spel genererar poäng med en hastighet av 5%; med följande undantag: Arabian Nights and Jackpottar 6000 genererar vid 5%; och Roulette, Blackjack,Jacks eller Better, Punto Banco, Baccarat, Casino Hold’em, Oasis Poker and TXS Hold’em genererar vid 1%. Klicka <a href="[Metadata:value(.FppRatesUrl)]">here</a> för en komplett lista över spel och deras priser.</li>
<li>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]förbehåller sig rätten att ändra eller avbryta
Cash Rewards erbjudande på bolagets eget gottfinnande.</li>
</ol>

