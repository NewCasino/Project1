Mitt sportkonto