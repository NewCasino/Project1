﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)]: r'Rollback Anmälan

