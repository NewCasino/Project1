Du kan inte göra en insättning.