﻿<p>Hej $FIRSTNAME$,</p>
<p>Ditt uttag har slutförts.</p>
<p>
  <span style="font-size: medium;">
    <strong style="color: #ff3366;">Kontrollera saldot på ditt bankkonto.</strong>
  </span>
</p>
<p>
  Tveka inte att kontakta oss om du har frågor. <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.
</p>
<p>
  Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet
</p>