Kina, Yuan Renminbi