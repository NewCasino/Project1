﻿/game/gamerules.jsp?game=blackjack2-3h&lang=sv