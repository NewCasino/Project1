﻿Betsoft spelande
