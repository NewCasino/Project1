﻿Annat
