Vänligen fyll i ditt lösenord