﻿/game/gamerules.jsp?game=tenhvideopokerdw&lang=sv