Vänligen välj din titel