﻿Vänligen ange ditt användarnamn
