﻿Uttag