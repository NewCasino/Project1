E-plånbok nummer