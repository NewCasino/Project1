﻿Typ