Ange bankens namn.