﻿Summa