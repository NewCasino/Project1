Mottagarens mobilnummer