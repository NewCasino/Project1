﻿Registrera ditt nya [Metadata:value(/Metadata/Settings.Operator_DisplayName)] konto 