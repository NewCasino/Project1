Skicka om verifieringskod ({0} sekunder)