﻿'linjär'