﻿Du måste välja en av de tillgängliga alternativen
