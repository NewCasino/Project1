﻿Emailfältet får inte lämnas tomt
