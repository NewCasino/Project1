Spelinformation