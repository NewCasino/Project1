﻿/game/gamerules.jsp?game=ice&lang=sv