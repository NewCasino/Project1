﻿Självexkludering till
