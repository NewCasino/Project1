﻿Inloggningen misslyckades. Du har valt att permanent självexkludera dig. Vill du ta bort din självexkludering, kommer du att få chansen att göra detta först efter ett år sedan du har självexkluderat dig.

