﻿Land Blockerad
