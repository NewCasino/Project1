﻿Går ut {0}
