﻿Oasis Poker Serier
