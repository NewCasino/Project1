﻿Misslyckades med att ladda saldo, var vänlig och prova igen senare.
