Vänligen ange din titel