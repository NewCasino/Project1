Uttag direkt till ditt NETELLER konto