﻿Visa menyn

