﻿Återstående omsättningskrav