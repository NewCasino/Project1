Kontakta oss