﻿Ny
