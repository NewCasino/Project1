Din e-post adress