Betala per telefon (Luxemburg)