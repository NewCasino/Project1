﻿({0} vinster totalt just nu)