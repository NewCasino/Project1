﻿Din adress måste innehålla minst två tecken
