Ange SMS-koden.