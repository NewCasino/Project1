Problem med casinots funktioner