﻿Använd standard
