Stäng