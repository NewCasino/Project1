﻿( frivilligt)


