﻿/game/gamerules.jsp?game=lrletitride2&lang=sv