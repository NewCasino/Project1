﻿Ditt innehåll här
