ID-nummer