Med E-pro kan du snabbt sätta in pengar från ditt kreditkort till ditt spelkonto. Ange bara dina kortuppgifter och så snart ditt kreditkort har verifierats kommer pengarna att föras över till ditt spelkonto, säkert och omedelbart.