﻿lottery
