Kreditera till {0} konto