Min favoritplats?