﻿Support
