﻿Roulette Pro Serier
