Kortägarens namn