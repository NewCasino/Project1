Ange ett mobilnummer med 7 till 30 siffror