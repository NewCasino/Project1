Uttag av pengar direkt till ditt SpeedCard-konto