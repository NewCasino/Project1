﻿De tillbakadragande transaktioner som anges nedan är närvarande.
Du kan avbryta dessa transaktioner och omedelbart återvända medel tillbaka till ditt konto genom att trycka rollback knappen.
Dina pengar kommer att finnas tillgängliga omedelbart på ditt konto.
