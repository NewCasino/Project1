Bekräfta lösenordet