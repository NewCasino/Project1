Utfärda en Ukash förbetald voucher och för över pengar till den nya vouchern.