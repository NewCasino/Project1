﻿När du klickar på ‘Bekräfta’, omdirigeras du direkt till Paykwik för att ange din voucherkod
