﻿UIPAS Konto-ID
