E-postadressens domän inte tillåten