﻿Bordsspel
