vecka