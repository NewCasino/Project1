Ange din kompis användarnamn.