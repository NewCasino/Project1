Glömt användarnamn