<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Syftet med detta e-mail är att bekräfta din lönegräns $LIMITAMOUNT$ $LIMITPERIOD$ kommer att tas bort den $LIMITEXPIRYDATE$. <br /><br /> Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p><br /> Vänliga Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kontaktsupport teamet</p>