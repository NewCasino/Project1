Uttag av pengar direkt till ditt eWire-konto