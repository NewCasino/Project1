Euteller är en direkt banköverföringsmetod online för finska banker.