﻿/game/gamerules.jsp?game=wizards&lang=sv