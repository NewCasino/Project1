﻿Betalare