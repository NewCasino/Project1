Kvitto