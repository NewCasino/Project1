﻿Fyll kontonummer