Beloppet överstiger din dagliga gräns