﻿Kampanjer
