﻿Sätt en sessionsgräns
