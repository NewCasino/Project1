﻿Bolivia