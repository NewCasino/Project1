Gör ett uttag direkt med ditt SpeedCard konto.