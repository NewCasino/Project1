﻿Uttag av pengar direkt till din bank via Alternative Payment Exchange