﻿Toppengaspelare
