Uttag direkt till ditt SOFORT konto