Kortnummer kan inte vara tomt.