Vänligen ange ditt Neteller Konto ID