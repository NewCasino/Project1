﻿Mobilprefix måste anges
