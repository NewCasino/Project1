﻿Självexkludering under 6 månader
