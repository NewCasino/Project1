<p>Du har begärt att din [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] e-mailadress ska ändras. En bekräftelse har skickats till den nya e-mail adressen($EMAIL$).</p><p>Om du inte har bet tom att ändra din e-mailadress, vänligen kontakta oss omedelbart på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p>Vänliga hälsningar, <br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>