Ange filialkoden.