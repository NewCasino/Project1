Verifieringskod kunde inte skickas, kontrollera ditt mobilnummer eller försök igen.