Du måste logga in för att kunna spela spelet.