﻿Gör ett uttag direkt till din bank via DengiOnline
