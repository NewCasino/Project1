Aktuella jackpots