Skapa ditt lösenord