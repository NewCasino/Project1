Valideringskoden består av 6 siffror.