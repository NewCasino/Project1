﻿/game/gamerules.jsp?game=bubbles&lang=sv