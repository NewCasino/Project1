Ange din adress