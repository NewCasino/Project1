Välj insättningskonto.