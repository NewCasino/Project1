Betala via SMS