﻿/game/gamerules.jsp?game=pandorasbox&lang=sv