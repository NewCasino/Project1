Total casino FPP poäng: