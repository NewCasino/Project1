Procentuell