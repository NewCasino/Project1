﻿Du spelar nu med riktiga pengar under jurisdiktionen i {0}.