﻿Fyll i onto holding filial