Veckovis gräns (var 7:e dag fr.o.m. tidpunkten då gränsen sattes)