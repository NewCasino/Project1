﻿Har du glömt ditt lösenord?
