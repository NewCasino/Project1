﻿DebitMisslyckades