Nyaste spelen