﻿/Kasino/FPP/Kurs
