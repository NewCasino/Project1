﻿Spelens RTP
