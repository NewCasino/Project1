﻿Bakåt
