Premie.