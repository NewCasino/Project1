﻿Double transaction request submit