﻿/game/gamerules.jsp?game=hrpuntobanco&lang=sv