﻿Sverige