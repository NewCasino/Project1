﻿Populära spel
