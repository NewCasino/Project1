Föreg<span class="Hideable">ious</span> {0} spel