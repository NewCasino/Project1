E-postadressen kan inte vara tom.