Spela {0} för riktiga pengar nu!