Återstående vadslagningskrav