﻿Skrivbord sidan
