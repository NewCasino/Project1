Insättning direkt till ditt Intercash kort