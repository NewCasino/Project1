﻿Endast nummer och komma är tillåtet. Vänligen använd punkt för decimalteckan och fyll i nummer utan formatering.
