Totalt antal jackpots