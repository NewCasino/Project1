Min favorithäst?