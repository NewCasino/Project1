﻿Jättipottipelit

