Misslyckades, kontrollera angivna uppgifter och försök igen.