Transaktionen kunde inte genomföras just nu.