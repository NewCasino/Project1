﻿Rabobank
