Födelsedatum