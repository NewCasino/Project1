﻿/game/gamerules.jsp?game=baccarat2&lang=sv