﻿Dölj Saldon
