﻿/game/gamerules.jsp?game=fortuneteller&lang=sv