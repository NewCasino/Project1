﻿Kasino Spel
