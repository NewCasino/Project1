Debet-voucherns kod