Kortnummer krävs