﻿<div class=" sitemap_items">
<div class="root_title">[Metadata:value(/Metadata/Settings.Operator_DisplayName)]</div>
<ul class=" items">
<li><a href="/">Hem</a></li>
<li><a href="/ help">Hjälp</a></li>
<li><a href="/customersupport">Kundsupport</a></li>
<li><a href="/deposit">Betalningsmetoder&nbsp;</a></li>
<li><a href="/ForgotPassword">Glömt Lösenord</a></li>
<li><a href="/register">Gå Med Nu</a></li>
<li><a href="#top">Logga in</a></li>
<li><a href="/Sports/Home ">Sport</a></li>
<li><a href="/Casino/Lobby">Casino</a></li>
<li><a href="/Poker/">Poker</a></li>
<li><a href="/Bingo/">Bingo</a></li>
<li><a href="/Promotions/Home">Kampanjer</a></li>
<li><a href="/AboutUs">Om Oss</a></li>
<li><a href="/ResponsibleGaming">Ansvarsfullt Spelande</a></li>
<li><a href=" /TermsConditions">Villkor &amp; </a></li>
<li><a href="/Sitemap">Webbkarta</a></li>
<li><a href="/Affiliate/Home">Dotterbolag</a></li>
</ul>
</div>
<div class="sitemap_items">
<div class="root_title">Sports</div>
<ul class="items">
<li><a href="/ help/Sports">FAQ</a></li>
<li><a href="/ Promotions/home/sportsbook">Kampanjer&nbsp;</a></li>
</ul>
</div>
<div class="sitemap_items">
<div class="root_title">Casino</div>
<ul class="items">
<li><a href="/help/Casino ">FAQ</a></li>
<li><a href="/Promotions/home/casino">Kampanjer</a></li>
</ul>
</div>
<div class="sitemap_items">
<div class="root_title">Poker</div>
<ul class="items">
<li><a href="#">Ladda ner klient</a></li>
<li><a href="/Poker/Tournaments/CAKEPoker">Turneringar</a></li>
<li><a href="/ PokerSchool">Poker Skola</a></li>
<li><a href="/ help/Poker">FAQ</a></li>
<li><a href="/ Promotions/TermsConditions/poker/LoyaltyLevels">LojalitetsNivåer</a></li>
<li><a href="/ Promotions/home/Poker">">Kampanjer</a></li>
</ul>
</div>
<div class=" sitemap_items">
<div class="root_title">Kampanjer</div>
<ul class="items">
<li><a href="/ Promotions/Home">Topp kampanjer</a></li>
<li><a href="/ Promotions/home/sportsbook">Sport</a></li>
<li><a href="/ Promotions/home/casino">Casino</a></li>
<li><a href="/ Promotions/home/Poker">Poker</a></li>
</ul>
</div>
<div class=" sitemap_items">
<div class=" root_title">Dotterbolag</div>
<ul class=" items">
<li><a href="/Affiliate/home">Logga in</a></li>
<li><a href="#">Glömt lösenordet??</a></li>
<li><a href="#">Registrera Dig Nu</a></li>
</ul>
</div>
