﻿<em>Det här meddelandet har skickats av en kund via sidan "Kontakta oss" på webbsidan.<br />
BESVARA INTE det här e-postmeddelandet direkt! Du hittar e-post för kundmeddelande nedan.</em>
<hr/>
<ul>
<li><strong>Kundens e-post</strong>:$EMAIL$</li>
<li><strong>Kundens namn</strong>:$NAME$</li>
<li><strong>Ämne</strong>:$SUBJECT$</li>
<li><strong>Användar-ID</strong>:$USERID$</li>
<li><strong>Användarnamn</strong>:$USERNAME$</li>
</ul>
<hr/>
<pre>$CONTENT$</pre>