Vänligen fyll i mottagarens telefonnummer. 