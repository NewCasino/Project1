﻿Överföring från dittr {0} konto