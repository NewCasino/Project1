Senaste kort