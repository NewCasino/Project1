Du har bara {0} poäng, vilket inte uppfyller minimikraven ({1} poäng).