﻿/game/gamerules.jsp?game=hrblackjackonedk&lang=sv