Godkänn