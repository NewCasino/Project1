﻿Alla turneringar
