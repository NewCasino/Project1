Om du är kvalificerad och har en bonuskod för en bonus, vänligen skriv den nedanför och tryck på skicka