Ja, skicka mig exklusiva erbjudanden via SMS. 