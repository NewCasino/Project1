﻿Stäng
