Min favoritsuperhjälte?