﻿Befintliga Kort
