﻿Endast nummer och komma är tillåtet. Vänligen använd punkt för decimaltecken och fyll i nummer utan formatering.
