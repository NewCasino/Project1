Debitera {0} konto.