﻿Ditt nya lösenord här
