﻿Videokolikkopelit

