Initialt omsättningskrav