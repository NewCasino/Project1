En permanent självuteslutningsperiod