Gammalt lösenord