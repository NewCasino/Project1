﻿Vänligen ange användarnamn och lösenord.


