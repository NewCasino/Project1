﻿Live Multispelare Roulette
