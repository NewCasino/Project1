Betala per telefon (Polen)