Uttag direkt till ditt ePay konto