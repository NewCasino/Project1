﻿Mobil betalning
