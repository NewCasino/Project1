﻿<!—Infoga Bakgrundsbild här -->

