Välj telefonnummerprefix