﻿Logga in

