﻿<img src="//cdn.everymatrix.com/_casino/2/272782A718C03124BC459616D30A5DBC.jpg" />
