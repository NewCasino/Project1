Betala per telefon (Spanien)