Hämta dina pengar