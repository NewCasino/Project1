﻿BANKLINKNORDEA