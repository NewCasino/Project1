﻿Visa Saldon
