Visa Delta/Debet