﻿/game/gamerules.jsp?game=lrblackjack2-3h&lang=sv