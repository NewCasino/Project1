Vänligen fyll i mottagarens mobilnummer