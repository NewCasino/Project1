Fel, det här spelet kan inte spelas i spela på skoj-läget!