Uttag av pengar direkt till ditt MasterCard.