﻿Bonusar
