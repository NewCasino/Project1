﻿Oddsbonus
