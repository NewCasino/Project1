Bonusbelopp