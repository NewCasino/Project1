﻿Uttag
