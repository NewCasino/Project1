﻿Klas Poker
