﻿Spela
