Visa populära bord