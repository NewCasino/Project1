casino FPP