Skicka nytt