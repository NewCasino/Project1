Sätt insättningsgräns