Visa alla kategorier