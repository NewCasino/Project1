﻿Ditt användarnamn här


