Smart SMS lösenord