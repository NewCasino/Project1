Filter - Betalningsalternativ