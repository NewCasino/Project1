Du kommer inte att kunna logga in på ditt bettingkonto under uteslutningsperioden på ett 1 år