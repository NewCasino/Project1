﻿/game/gamerules.jsp?game=jacksorbetter10&lang=sv