Överför pengar via {0}