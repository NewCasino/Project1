Vänligen välj datum giltigt från