Bankkontonr.