Ange NIP.