﻿Odds Bonus
