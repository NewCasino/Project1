﻿/game/gamerules.jsp?game=shvideopokerjob&lang=sv