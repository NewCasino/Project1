Sverige, Kronor