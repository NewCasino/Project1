﻿Validation kod