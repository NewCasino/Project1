Vinnare nu