﻿You have requested an amount above {$}. Please try again.