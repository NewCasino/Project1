Du kommer inte att kunna logga in på ditt konto under den valda tidsperioden.