Självavstängning