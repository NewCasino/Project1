Visa spel i standardordning