﻿€ (EUR)