Aktivera bakgrunden