﻿Utbetala
