Transaktionen är inte slutförd.