﻿{0}

