﻿{0}t sedan