﻿<p>Hej $FIRSTNAME$,</p>
<p>Din insättning lyckades.</p>
<p>
  <span style="font-size: medium;">
    <strong style="color: #ff3366;">Klicka på knappen "Uppdatera" (INTE uppdateringsknappen på webbläsaren) överst på sidan för att ladda om saldot.</strong>
  </span>
</p>
<p>
  Tveka inte att kontakta oss om du har frågor. <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.
</p>
<p>
  Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet
</p>