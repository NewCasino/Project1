﻿Avslutas vid {0}
