﻿Referens-ID