﻿Source and destination accounts are the same