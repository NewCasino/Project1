Ladda fler spel nu!