﻿[Metadata:value(/Metadata/GammingAccount/CakeNetwork.Display_Name)] Kredit & Debet

