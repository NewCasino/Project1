﻿Fel UIPAS Konto-ID
