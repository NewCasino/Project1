Stänger kl.