Biljettpris