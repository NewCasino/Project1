Transaktionen har avbrutits.