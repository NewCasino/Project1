﻿/game/gamerules.jsp?game=pacific&lang=sv