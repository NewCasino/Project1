Ange ditt postnummer