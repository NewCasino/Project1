﻿...eller