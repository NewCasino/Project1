Du måste vara äldre än {0} år