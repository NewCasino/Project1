Ange sessionsgräns