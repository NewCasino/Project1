﻿Insättning med TLNakit
