﻿Generera Kod
