﻿Avsluta
