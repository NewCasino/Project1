﻿/game/gamerules.jsp?game=mansion&lang=sv