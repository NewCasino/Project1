﻿Spelande
