﻿Logga in på din onlinebank för att fullfölja betalningen
