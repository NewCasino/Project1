﻿Your request could not be completed. Please call NETELLER Customer Service.