Skicka verifieringskod