﻿Din bonuskod
