Qiwi är en eWallet och terminalservice som erbjuder dig säkra betalningsmetoder. 