﻿Netherlands Antilles