En 3-månaders självuteslutningsperiod