E-postadressen verkar felstavad.