<div id="help-area">
    <h3 class="content-item" id="1">
        <strong>Allmänna regler</strong>
    </h3>
    <ol class="ord-list">
        <li>Alla insatser godkända av [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; omfattas av dessa regler.</li>
        <li>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; förbehåller sig rätten att annullera insatser som görs på uppenbart "dåliga" odds, ändrade odds eller en insats som görs efter att en tävling startat.</li>
        <li>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; förbehåller sig rätten att vägra, insränka, annullera eller begränsa en insats.  </li>
        <li>Satsningar graderas först när tävlingen avgjorts.</li>
        <li>Vinnaren av en tävling kommer att fastställas det datum då tävlingen avgörs, [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; erkänner inte protest- eller upphävda beslut för insatser. Resultat för en tävling som avbryts efter starten av tävlingen kommer att beslutas mot bakgrund av reglerna som anges för denna idrott genom [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp;.</li>
        <li>Enligt lagarna för the Lottery and Gaming Authorities in Malta har ingen under 18 år tillstånd att göra en insats.</li>
        <li>Alla regler, föreskrifter och satsningar häri är föremål för ändringar och revideringar av [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; utan föregående skriftligt meddelande.</li>
        <li>Maximalt insatsbelopp på alla idrottsevenemang kommer att fastställas genom [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; och kan ändras utan föregående skriftligt meddelande. [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; förbehåller sig också rätten att justera gränserna för individuella konton.</li>
        <li>I de fall pengar krediteras till ett kundkonto av misstag åligger det kunden att underrätta [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; om ovannämnda fel utan dröjsmål. För konton med minussaldo, förbehåller sig [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; rätten att annullera alla pågående spel, oavsett om placerats med medel till följd av fel eller inte.</li>
        <li>Medlemmar är själva ansvariga för sina kontotranskationer. Se till att granska och bekräfta dina insatser för eventuella fel innan du skickar in dem. När en transaktion är klar, kan den inte ändras. [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; tar inte ansvar för försvunna eller duplicerade satsningar som görs av kunden och kommer inte att ta under övervägande begäran om differens därför att ett spel saknas eller dupliceras. Kunder granska sina transaktioner i "Mitt Sports Betting konto" på webbplatsen efter varje session för att garantera att alla begärda satsningar godtogs.</li>
        <li>Tvister skall göras inom sju (7) dagar från den dag insatsen i fråga har beslutats. Inga krav kommer att godtas efter denna tidsfrist. Kunden är ensamt ansvarig för sina kontotransaktioner.</li>
        <li>Alla saldon och transaktioner visas i den valuta markerad när kontot ursprungligen öppnades.</li>
        <li>Vinster kommer alltid att beräknas med hjälp av European Odds. Observera att när du konverterar odds till brittisk standard, kan avrundningsfel förekomma, då vissa odds inte har en exakt översättning till bråk i brittisk stil. Här kommer vi att visa närmaste bråkodds.</li>
        <li>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; förbehåller sig rätten att stänga ett kundkonto utan uppsägningstid och returnera alla medel till vederbörandes huvudsakliga plånbok.</li>
        <li>I händelse av en diskrepans mellan den engelska versionen av dessa regler och alla andra språk, kommer den engelska versionen att anses vara korrekt.</li>
        <li>Ackumulatorer (Parlays, Multis): Vi tar emot upp till 10 resultat i en ackumulator. Om vissa resultat är "ömsesidigt beroende", exempel: placera insats på Chelsea för att vinna engelska Premier League kombinerat med en hemmavinst i det sista avgörande spelet, kommer dessa insatser vara ogiltiga. </li>
    </ol>
    <h3 class="content-item" id="2">
        <strong>Fotboll</strong>
    </h3>
    <ol class="ord-list">
        <li class="content-statement">
            <strong>Kommer spelaren göra mål</strong>: Ingen återbetalning på icke startande
        </li>
        <li class="content-statement">
            <strong>Förste Målskytt</strong>: Ingen återbetalning på icke startande
        </li>
        <li class="content-statement">
            <strong>Sista Målskytt</strong>: Ingen återbetalning på icke startande
        </li>
        <li class="content-statement">
            <strong>Första Lag att göra Mål</strong>:
        </li>
        <li class="content-statement">
            <strong>Tidpunkt för Första Mål</strong>: Bets are settled on what time the goal is actually scored from official source
        </li>
        <li class="content-statement">
            <strong>Last Team to score</strong>: In the event of an abandoned game bets stand on scores that have taken place already, Extra Time does not count for these markets.
        </li>
        <li class="content-statement">
            <strong>Race To X Goals</strong>: Settled on the team who reaches the quoted number of goals first in the event of an abandonment before 90 minutes have been played then all bets will be void unless settlement is already determined.
        </li>
        <li class="content-statement">
            <strong>Both Team To Score</strong>: Baserat på om bägge lagen gör mål i matchen.
        </li>
        <li class="content-statement">
            <strong>Team Score Over Under</strong>: Based on total number of goals scored by a team in the match. Extra Time goals are not included.
        </li>
        <li class="content-statement">
            <strong>Antal mål</strong>: Spel på Antalet Mål inkluderar "egna mål"
        </li>
        <li class="content-statement">
            <strong>Goal In Time Range</strong>: Will be the official time of goal scored that will count. Extra Time not included
        </li>
        <li class="content-statement">
            <strong>Att Göra Mål I Båda Halvlekarna</strong>: Is a Yes/No Bet if a Team/Teams will score in both halves.
        </li>
        <li class="content-statement">
            <strong>To Win To Nil</strong>: Team to win the match and keep a clean sheet.
        </li>
        <li class="content-statement">
            <strong>Vinstmarginal</strong>: Settled on the result of game. The teams will be given various margins of winning and it will be the final result that counts.
        </li>
        <li class="content-statement">
            <strong>To Win Either Half</strong>: A Team needs to win minimum one of the two halves in order for this bet to winning.
        </li>
        <li class="content-statement">
            <strong>To Win Both Halves</strong>: The team must score more goals than the opposition in both halves of the match.
        </li>
        <li class="content-statement">
            <strong>Komma Från Underläge Och Vinna</strong>: Laget måste ligga under i någon fas av matchen, men till slut vinna matchen i 90 minuter fulltid.
        </li>
        <li class="content-statement">
            <strong>Corners Over Under</strong>: Based on a specific line added in Over/Under for corners taken in the match. Extra Time does not count
        </li>
        <li class="content-statement">
            <strong>Antal hörnor</strong>: Baserat på totala antalet hörnor tagna i matchen.
        </li>
        <li class="content-statement">
            <strong>Vem Gör Först X Hörnor</strong>: Settled on the team who reach the quoted number of corners first, in the event of an abandonment before 90 minutes have been played then all bets will be void unless settlement is already determined.
        </li>
        <li class="content-statement">
            <strong>Tid För Nästa LagMål</strong>: Settlement will be made by the time given by the official match source as the time of First/Next goal is scored.
        </li>
        <li class="content-statement">
            <strong>Varningar Över/Under</strong>:
        </li>
        <li class="content-statement">
            <strong>Lag Varningar Över/Under</strong>: Settlement will be made with reference to all available evidence to cards shown during the scheduled 90 minutes play. Any card shown after the full time whistle has been blown will be disregarded.
        </li>
        <li class="content-statement">
            <strong>Half With Most Corners</strong>: According to the corner numbers of each half, the half with more corners won
        </li>
        <li class="content-statement">
            <strong>Lag Antal Hörnor</strong>: Number of corners a team gets
        </li>
        <li class="content-statement">
            <strong>Last Corner Kick</strong>: Which team will get the last corner kick, based on the current corner
        </li>
        <li class="content-statement">
            <strong>Clean Sheet</strong>: Team who keeps a clean sheet won
        </li>
        <li class="content-statement">
            <strong>Most Corners</strong>: Team that gets more corners in a match will win
        </li>
        <li class="content-statement">
            <strong>Nästa hörna</strong>: Which team will get the next corner, based on the current corner
        </li>
        <li class="content-statement">
            <strong>MatchSpel Och Totaler</strong>: Combine 1x2 and over under, only both won bets will win, all others lost
        </li>
        <li class="content-statement">
            <strong>Att Gå Till övertid</strong>: If match goes to overtime, then won, if  not, lost
        </li>
        <li class="content-statement">
            <strong>Utvisning</strong>: Will there be red cards or not
        </li>
        <li class="content-statement">
            <strong>Hörnor Udda/Jämt</strong>: Total corners are Odd or Even
        </li>
        <li class="content-statement">
            <strong>LagMål Inom Tidsintervallet</strong>: Will be the official time of goal scored that will count. Extra Time not included
        </li>
        <li class="content-statement">
            <strong>Lag Hörnor Udda/Jämt</strong>: Team total corners are odd or even
        </li>
        <li class="content-statement">
            <strong>Lag Hörnor Över/Under</strong>: Team total corners over or under a parameter
        </li>
        <li class="content-statement">
            <strong>Att Gå Till Straffar</strong>: Will the match go to penalty time?
        </li>
        <li class="content-statement">
            <strong>En Inbytare Att Göra Mål</strong>: Will a substitute score a goal
        </li>
        <li class="content-statement">
            <strong>Antal Kort</strong>: Settlement will be made with reference to all available evidence to cards shown during the scheduled 90 minutes play. Any card shown after the full time whistle has been blown will be disregarded.
        </li>
        <li class="content-statement">
            <strong>Gula Kort Udda/Jämt</strong>: Settlement will be made with reference to all available evidence to cards shown during the scheduled 90 minutes play. Any card shown after the full time whistle has been blown will be disregarded.
        </li>
        <li class="content-statement">
            <strong>Första Lag Varning</strong>: Which team will get the next card, accordingly to the current card
        </li>
        <li class="content-statement">
            <strong>SjälvMål Görs</strong>: Will there be own goal scored?
        </li>
        <li class="content-statement">
            <strong>Metod För Vinst</strong>: How the match ends to get a winner
        </li>
        <li class="content-statement">
            <strong>Lag Att Erhålla Det Första Gula Kortet</strong>: Which team to receive the next yellow card, according to the current card
        </li>
        <li class="content-statement">
            <strong>Högsta Antal Mål Under Halvlek</strong>: Half with most goal wins
        </li>
    </ol>

    <h3 class="content-item" id="3">
        <strong>Tennis</strong>
    </h3>
    <ol class="ord-list">
        <li class="content-statement">In case of retirement, disqualification or change of surface mid-match, all bet's which cannot be settled by current score will be voided</li>
        <li class="content-statement">(1) A set is abandoned at 4-4: bets on Over/Under 7.5 games or fewer in the set are settled as winners/losers respectively; bets on ex Over/Under 10.5 games or more are void.</li>
        <li class="content-statement">Sets Betting: If a tennis match is not completed because of a player retirement or disqualification, all not decided set bets will be considered void.</li>
        <li class="content-statement">Delay or Suspension: If a tennis match is completed, all bets stand as written. A delay in the start of a match will not affect the standing of bets, nor will a suspension, as long as play is resumed and the match completed;</li>
        <li class="content-statement">In the event a match does not go the specified number of sets, and the match is shortened by tournament officials, the leader determined to be official by tournament officials shall be the winner;</li>
        <li class="content-statement">Example: A match is scheduled for 5 sets, but only 3 sets can be played because of weather. The leader at the end of 3 sets would be declared the winner of the match.</li>
        <li class="content-statement">
            <strong>Tie Break</strong>: If there is tie break, won, if no, lost
        </li>
        <li class="content-statement">
            <strong>Game Score</strong>: Exact score of the game and will the server be broken
        </li>
        <li class="content-statement">
            <strong>Game To Deuce</strong>: Will there be 40:40 in a game?
        </li>
        <li class="content-statement">
            <strong>Games Won Over Under</strong>: Total games of a player are over or under a parameter
        </li>
        <li class="content-statement">
            <strong>Antal Spelade</strong>: Total games of both players in a set
        </li>
        <li class="content-statement">
            <strong>Att Vinna Åtminstonde Ett Set</strong>: If a player wins 1 set or not when the match ends
        </li>
        <li class="content-statement">
            <strong>Race To X Games</strong>: Who will win the x game in x set
        </li>
        <li class="content-statement">
            <strong>Vem Gör Först X Poäng</strong>: Which player will win xth point, game y, n set
        </li>
        <li class="content-statement">
            <strong>Poäng handicap</strong>: Who will win the game with the handicap parameter in that set
        </li>
        <li class="content-statement">
            <strong>Points Over Under</strong>: Total game points over under in x game, n set
        </li>
        <li class="content-statement">
            <strong>Points Won Over Under</strong>: Total points by each player, in x game, n set
        </li>
        <li class="content-statement">
            <strong>To hold first service game</strong>: Will the player hold the first service game in first set?
        </li>
        <li class="content-statement">
            <strong>Game Of First Service Break</strong>: First service break is in which game at first set
        </li>
        <li class="content-statement">
            <strong>Total Service Breaks</strong>: How many service breaks will be in 1st set
        </li>
        <li class="content-statement">
            <strong>Vinstmarginal</strong>: What is the difference of total number of games won by winner and loser
        </li>
        <li class="content-statement">
            <strong>Lose 1st Set And Win The Match</strong>: Which player lost 1st set but won the match in the end
        </li>
    </ol>

    <h3 class="content-item" id="4">
        <strong>Amerikansk fotboll, rugby och AFL</strong>
    </h3>
    <ol class="ord-list">
        <li>Minsta tid för gällande: När det gäller insatser, fastställs vinnare och förlorare av slutresultatet (inklusive övertid), förutsatt att matchen pågått i minst 55 minuter.</li>
        <li>Om en match avbryts efter 55 minuter och inte återupptas samma dag, kommer oavsett om matchen avslutas vid en senare tidpunkt, kommer poängen när spelet stoppas att avgöra insats resultatet.</li>
        <li>Om matchen avbryts före slutförandet av 55 minuter och inte återupptas samma dag, kommer alla insatser noteras som "inte gällande" och pengarna återbetalas.</li>
        <li>Alla insatser på matchen kommer att inkludera övertidsmål om inte annat anges.</li>
        <li>Om inte känt före en tävling, måste alla tävlingar spelas på planerat datum och på det planerade området för att gälla.</li>
        <li>Australian Rules, Rugby League, Super League och Rugby Union. Insatser kommer att betalas på det slutliga resultatet för en tävling (normaltid eller extratid i förekommande fall).</li>
        <li>NFL Propositioner rangordnas genom att använda resultaten som anges på www.NFL.com.</li>
        <li>Arena Football Propositioner rangordnas genom att använda resultaten som anges på www.Arenafootball.com.</li>
    </ol>
    <h3 class="content-item" id="5">
        <strong>Ishockey</strong>
    </h3>
    <ol class="ord-list">
        <li>Om inget annat anges, gäller insatser ENDAST för ordinarie tid och inkluderar inte heller övertid eller straffsparkar. Exempel: Det står 3-3 mellan Rangers och Kings efter ordinarie tid och går vidare till övertid. Rangers vinner till slut. Slutresultat för insats är Rangers 3, Kings 3.</li>
        <li>Om en rad inkluderar övertid, ska det tydligt anges i spelerbjudandet och vara tydligt skrivet på biljetten. Kontrollera din biljett noggrant.</li>
        <li>Straffsparkar är uttryckligen en del av övertid. Vid straffsparkar krediteras vinnaren med ett extra mål.</li>
        <li>Exempel: Det står 2-3 mellan Dynamo och CSKA och går vidare till straffsparkar. Dynamo vinner straffarna, För vår radmatch "Dynamo inklusive OT" vs. "CSKA inklusive OT", slutresultatet för insats är Dynamo 3, CSKA 2.</li>
        <li>Minsta tid för Action: Matcher måste spelas minst 55 minuter för att gälla. Om en match avbryts innan 55 kompletta minuter har spelats, lämnas alla insatser på resultatet av matchen tillbaka.</li>
    </ol>
    <h3 class="content-item" id="6">
        <strong>Handboll</strong>
    </h3>
    <ol class="ord-list">
        <li>För insatser, avgörs vinnare och förlorare av ställningen vid ordinarie tids utgång. Extratid (en förlängning av ordinarie tid) kommer inte att räknas om inte annat anges.</li>
        <li>Om en match blir uppskjuten av någon anledning, kommer alla insatser att annulleras och pengarna betalas tillbaka om matchen inte schemaläggs att spelas inom 24 timmar efter den ursprungliga tiden för avspark.</li>
        <li>Om en matcharena ändras kommer redan placerade insatser gälla förutsatt att hemmalaget fortfarande är angivet. Om hemma- och bortalaget för en registrerad match ändras kommer insatser placerade på  den ursprungliga registreringen att vara ogiltiga.</li>
        <li>
            Game props: Alla game props, inklusive följande aktiviteter, kommer uteslutande att avgöras på ordinarie tid och exkludera eventuell övertid:
            <ol type="disc">
                <li>Spelresultat ojämn/jämn</li>
                <li>Dubbla resultat</li>
            </ol>
        </li>
    </ol>
    <h3 class="content-item" id="7">
        <strong>Basketball</strong>
    </h3>
    <ol class="ord-list">
        <li>Minsta tid för gällande: NBA-matcher måste spelas minst 43 minuter för att gälla. För alla andra basketligor, måste matcher spelas i minst 35 minuter om inte annat anges.</li>
        <li>När det gäller insatser, fastställs vinnare och förlorare av slutresultatet (inklusive övertid), förutsatt att spelet pågått den minsta tid som anges ovan. Om en match avbryts efter den minsta tiden har spelats och inte återupptas samma dag, kommer oavsett om matchen avslutas vid en senare tidpunkt, poängen när spelet stoppas att avgöra insats resultatet.</li>
        <li>Om spelet avbryts före den minsta tiden har uppnåtts och inte återupptas samma dag, kommer alla insatser noteras som "inte gällande" och pengarna återbetalas.</li>
        <li>Alla insatser på spelet kommer att inkludera övertidsmål om inte annat anges.</li>
        <li>Om inte känt före en tävling, måste alla tävlingar spelas på planerat datum och på den planerade platsen för att gälla.</li>
        <li>Dessa regler gäller både collage och profesionell basket.</li>
        <li>NBA resultat graderas med hjälp av statistik från NBA.com.</li>
        <li>NCAA Basketball resultat graderas med hjälp av statistik från espn.com.</li>
        <li class="content-statement">
            <strong>Dubbelchans</strong>: What will be the match result, double the result, 12, 1X, 2X
        </li>
        <li class="content-statement">
            <strong>Högsta Antal Mål Under Quarter</strong>: Quarter total points, highest quarter won
        </li>
        <li class="content-statement">
            <strong>Att Gå Till övertid</strong>: Will the match have Overtime play?
        </li>
        <li class="content-statement">
            <strong>Vem Gör Först X Poäng</strong>: Which team will win xth point
        </li>
        <li class="content-statement">
            <strong>Vinstmarginal</strong>: The margin between two teams, how many points will a team won
        </li>
        <li class="content-statement">
            <strong>Team Score Over Under</strong>: Total points of a team over or under a parameter
        </li>
        <li class="content-statement">
            <strong>Lag Udda/Jämt</strong>: Total points of a team are odd or even
        </li>
        <li class="content-statement">
            <strong>Last Team to score</strong>: Which team will get the last score based on the current scores
        </li>
        <li class="content-statement">
            <strong>Första Lag att göra Mål</strong>: Which team will score first
        </li>
        <li class="content-statement">
            <strong>Halvtid/Fulltid</strong>: Who will win first half and the match
        </li>
        <li class="content-statement">
            <strong>Högsta Antal Mål Under Halvlek</strong>: Half with most goal wins
        </li>
        <li class="content-statement">
            <strong>Which team wins jump ball</strong>: Which  team will have the first  possession/jumpball
        </li>
        <li class="content-statement">
            <strong>Points Won Over Under</strong>: Total points of a player is over or under a parameter
        </li>
        <li class="content-statement">
            <strong>Point Winner</strong>: Which player will get the xth point
        </li>
    </ol>

    <h3 class="content-item" id="8">
        <strong>Baseboll</strong>
    </h3>
    <ol class="ord-list">
        <li>När man satsar på antal totalt antal varv (over/under) måste matchen spelas i 9 omgångar (8.5 om hemmalaget leder) för att gälla. Om en match dömer eller suspenderar in extra omgångar, kommer resultatet avgöras efter den sista fulla omgången om inte hemmalaget gör oavgjort, eller tar ledningen i den nedre halvan av omgången, i vilket fall poängen avgörs när matchen döms.</li>
        <li>Resultatet för en match är officiell efter 5 omgångars spel om inte hemmalagat leder efter  4.5 omgångar. Om en match dömer eller suspenderar in extra omgångar, kommer vinnaren avgöras enligt den sista fulla omgången om inte hemmalaget gör oavgjort, eller tar ledningen i den nedre halvan av omgången, i vilket fall vinnaren avgörs när matchen döms. Alla pengar kommer att betalas tillbaka om hemmalaget gör oavgjort och sedan avbryts.</li>
        <li>[Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; godkänner inte uppskjutna spel, protester eller upphävda beslut om insatser. Alla insatser på baseball ska göras den angivna dagen, för att det ska gälla annars betalas alla pengar tillbaka.</li>
        <li>Money-line insatser på baseboll kommer att godkännas som gällande oavsett start-pitcher.</li>
        <li>MLB farmarligor: Om en dubbelmatch spelas mellan Lag A och Lag B och [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; sätter ett pris för Lag A vs. Lag B för endast en match, utan att beteckna det som antingen Spel 1 eller Spel 2, ska priset avse match 1. Om, i själva verket, Match 1 redan har startat, ska det avse Match 2.</li>
        <li>MLB Prop Rules: För prop, måste spelet gå 9 omgångar (8.5 om hemmalaget leder) för att gälla.</li>
        <li>MLB Propositioner rangordnas genom att använda resultaten som anges på www.MLB.com.</li>
    </ol>
    <h3 class="content-item" id="9">
        <strong>Volleyball</strong>
    </h3>
    <ol class="ord-list">
        <li>Om en match avbryts innan full tid uppnås och inte avslutas samma dag, betraktas insatser på matchresultat som ogiltiga och alla insatser skall återlämnas.</li>
        <li>Byte av arena: Om en matcharena ändras kommer redan placerade insatser gälla förutsatt att hemmalaget fortfarande är angivet. Om hemma- och bortalaget för en registrerad match ändras kommer insatser placerade på  den ursprungliga registreringen att vara ogiltiga.</li>
    </ol>
    <h3 class="content-item" id="10">
        <strong>Snooker</strong>
    </h3>
    <ol class="ord-list">
        <li>Match-up insats är baserat på korrekt markera den spelare som officiellt vinner matchen. Om en match startar &ndash; med servegenombrott för den första bilden &ndash; men av någon anledning inte avslutas, kommer den spelare som fortsätter till nästa omgång (eller förklaras vinnare av tävlingen/mästerskapet) att betraktas som vinnare. Skulle en match inte starta, kommer alla insatser att betalas tillbaka.</li>
        <li>Frame betting baseras på att korrekt markera slutresultatet för en snookermatch. I händelse en match startar men inte avslutas av någon anledning eller att en match inte startar, betalas alla insatser tillbaka.</li>
    </ol>
    <h3 class="content-item" id="11">
        <strong>Fighting</strong>
    </h3>
    <ol class="ord-list">
        <li>När klockan ljuder för att starta den första omgången kommer figthen anses vara officiell för insatser, oavsett om den planerade längden eller titel.</li>
        <li>En fight är en Technical Draw när en fight avslutas före ett anvisat antal omgångar. Detta är vanligtvis på grund av en oavsiktlig head-butt eller foul.</li>
        <li>En fight som betraktas som "ingen tävling" kommer att betala tillbaka alla insatser.</li>
        <li>Om insatsen erbjuden på en match omfattar draw som ett tredje alternativ och matchen slutar oavgjort, kommer satsningar på oavgjort betalas ut, kommer satsningar på båda de båda tävlande att gå förlorade. Om insatserbjudandet endast inkluderar de två boxarna, med oavgjort antingen inte erbjuds eller erbjuds som ett separat förslag, och matchen slutar oavgjort, kommer satsningar på endera boxaren återbetalas.</li>
        <li>En Over/Under (totalt) registrerad på en fight representerar det total antalet genomförda omgångar. Halvtid i en omgång är exakt en minut och trettio sekunder in i en treminuters omgång. Därmed skulle 9 ½ omgångar vara en minut och trettio sekunder av den 10:e omgången. Halvtid i en tvåminuters omgång är exakt en minut. Halvtid i en femminuters omgång är två och en halvminut.</li>
        <li>Resultaten kommer att graderas på grundval av det officiella resultatet vid boxningsringen. Resultaten är inte officiell för satsningar förrän de har kontrollerats av funktionärer vid boxningsarenan. Officiella eller inofficiella påföljder rörande ett beslut om en fight på grundval av överklagande, rättsprocess, rättegången, drogtestresultat, eller någon annan påföljd kommer godkännas för satsningar.</li>
        <li>Om inte annat anges måste matchen gå inom trettio dagar efter det planerade datumet för att insatser ska gälla.</li>
    </ol>
    <h3 class="content-item" id="12">
        <strong>Bandy</strong>
    </h3>
    <ol class="ord-list">
        <li>Om inget annat anges, är alla insatser endast för ordinarie tid och inkluderar inte heller övertid. I turneringar om en ny aktivetet formas i slutet av ordinarie tid, t ex vinna på övertid, då gäller straffsparkar.</li>
        <li>Speltid: Om formatet på en match ändras oavsett skäl från 2 x 45 minuter till 3 x 30 minuter, gäller alla satsningar utom insatser som hänvisar till antingen första eller andra halvlek.</li>
        <li>Byte av arena:Om en matcharena ändras kommer redan placerade insatser gälla förutsatt att hemmalaget fortfarande är angivet. Om hemma- och bortalaget för en registrerad match ändras kommer insatser placerade på den ursprungliga registreringen att vara ogiltiga.</li>
    </ol>
    <h3 class="content-item" id="13">
        <strong>Innebandy</strong>
    </h3>
    <ol class="ord-list">
        <li>För insatser, avgörs vinnare och förlorare av ställningen vid ordinarie tids utgång. Förlängning eller sudden death räknas inte med mindre än att så anges.</li>
        <li>Om en match avbryts innan full tid uppnås och inte avslutas samma dag, betraktas insatser på matchresultat som ogiltiga och alla insatser skall återlämnas.</li>
        <li>Om en match blir uppskjuten av någon anledning, kommer alla insatser att annulleas och alla insatser återbetalas.</li>
    </ol>
    <h3 class="content-item" id="14">
        <strong>Pilkastning</strong>
    </h3>
    <ol class="ord-list">
        <li>Insats på match: Den spelare som går vidare till nästa omgång kommer att betraktas som vinnare, förutsatt att en av spelarna kastat en pil i början av den första omgången. Om den första pilen inte kastas, kommer alla insatser att annulleras.</li>
        <li>Insats på set: Det totala antalet set som krävs för att vinna matchen måste fullföljas. Om av någon anledning matchen tilldelas någon av deltagarna innan det fulla antalet set är klart, annulleras alla insatser.</li>
    </ol>
    <h3 class="content-item" id="15">
        <strong>Futsal</strong>
    </h3>
    <ol class="ord-list">
        <li>Om inte annat anges, avgörs alla insatser endast på ordinarie tid. Detta omfattar två perioder av spel och den tid domaren lägger till som kompensation för skador och andra avbrott. Det inkluderar inte perioder av övertid eller straffsparkar.</li>
        <li>Om en match avbryts innan full tid uppnås och inte avslutas samma dag, betraktas insatser på matchresultat som ogiltiga och alla insatser skall återlämnas.</li>
        <li>Startdatum och tider för futsal som visas på vår webbsida är en indikation och kan inte garanteras vara korrekt. Om en match blir uppskjuten, kommer alla insatser gälla 48 timmar efter avspark. Om vi får information att en uppskjuten match har lagts till en tid efter två dagar kommer vi omedelbart lämna tillbaka alla medel från pågående satsningar.</li>
        <li>Byte av arena: Om en officiell ändring av arena sker efter det att insatser gjorts kommer dessa insatser att annulleras.</li>
    </ol>
    <h3 class="content-item" id="16">
        <strong>Poker</strong>
    </h3>
    <ol class="ord-list">
        <li>Spelare som placeras det högsta beloppet pengar kommer att vinna.</li>
        <li>För direkta insatser, måste tävlande starta i tävlingen för att de ska gälla.</li>
    </ol>
    <h3 class="content-item" id="17">
        <strong>Curling</strong>
    </h3>
    <ol class="ord-list">
        <li>Om inte annat anges ingår alltid extra ends alltid resultatet för insatser.</li>
        <li>För att en insats ska gälla, måste minst 6 ends fullföljas.</li>
        <li>Slutresultatet för en match är den poäng som rapporteras av turneringsorganisatörer. [Metadata:value(/Metadata/Settings.Operator_DisplayName)]&nbsp; respekterar varje turnerings poängregler och regler avseende godkända matcher.</li>
        <li>Insatser på matcher som skjuts upp eller suspenderas av någon anledning (till exempel, men inte begränsats till: Försämrade isförhållanden, elavbrott, eller schemaläggningsproblem) betraktas som "gällande" och kommer att graderas när turneringsorganisatörerna förkunnar att matchen avslutats.</li>
    </ol>
    <h3 class="content-item" id="18">
        <strong>Bordtennis</strong>
    </h3>
    <ol class="ord-list">
        <li>I händelse att en match startar men inte slutförs av någon anledning kommer alla insatser på resultatet av matchen betraktas som ogiltigt.</li>
        <li>Insats på set (Korrekt poäng) hänvisar till korrekt slutresultat i set.</li>
        <li>När det gäller lagmatcher, i händelse att en matchup mellan spelare spelas två gånger, gäller endast det första resultatet.</li>
    </ol>
    <h3 class="content-item" id="19">
        <strong>Galoppsport</strong>
    </h3>
    <ol class="ord-list">
        <li class="no-bullet">
            <h4>General</h4>
            <ol>
                <li class="help-li">All bets are settled in accordance with the official result at the time of the "weigh in". Any change to a result after this point will not count;</li>
                <li class="help-li">Walkovers and void races count as races but any horse involved will be treated as a non-runner.</li>
            </ol>
            <h4>Non-Runners och avhopp</h4>
            <ol>
                <li class="help-li">If a horse is withdrawn before coming under starter's orders, or is officially deemed by the starter to have taken no part in the race, then all bets on that horse are void. Your stakes will be returned on the withdrawn horse.</li>
            </ol>
            <h4>Non-Runners och avhopp</h4>
            <h4>Tidigt på morgonen priser/priser för tävlingar samma dag</h4>
            <ol>
                <li class="help-li">After the final declarations stage, Non-Runner no-bet will apply.</li>
            </ol>
            <h4>Dubbla uppdrag</h4>
            <ol>
                <li class="help-li">Where a horse is doubly engaged (named as a runner in more than one race) the bet will stand as a bet for the timed race. If the selection runs in the other race it would be treated as a non runner.</li>
            </ol>
            <h4>Re-runs</h4>
            <ol>
                <li class="help-li">In the event of a false start or any other incident resulting in a race being re-run, 'under starter's orders' is negated and stakes will be refunded on horses taking no part in the re-run;</li>
            </ol>
            <h4>Uppskjutanden</h4>
            <ol>
                <li class="help-li">If a race is abandoned or declared void then any bets will be void. If the race is postponed to a future day and the final Declarations stand, all bets will stand;</li>
                <li class="help-li">
                    However, all single bets on horse racing will be made void and any selection involved in accumulative bets will be treated as a non-runner if:
                    <ol>
                        <li class="help-li">The race is abandoned;</li>
                        <li class="help-li">The race is officially declared void;</li>
                        <li class="help-li">The conditions of the race are altered after bets have been made;</li>
                        <li class="help-li">The venue is altered;</li>
                        <li class="help-li">The running surface is altered (e.g. from Turf to All Weather).</li>
                    </ol>
                </li>
            </ol>
            <h4></h4>
            <h4>Ante-Post Betting</h4>
            <ol>
                <li class="help-li">Ante post betting will cease at the Final Declaration stage and all bets after this will be non-runner, no bet ;</li>
                <li class="help-li">Unless specifically stated otherwise, stakes are lost on an Ante-Post bet if a horse does not take part. </li>
                <li class="help-li">On days when classic or other trials occur, Ante-Post betting may be suspended and new prices issued;</li>
                <li class="help-li">Ante-Post bets on horses compulsorily withdrawn will be void and stakes returned. (Stewards are empowered to reduce the numbers in a race if, at the overnight declaration stage, too many have been left in for the safety of horses and jockeys. Jockey Club Rule 121). </li>
                <li class="help-li">Ante-Post bets are settled at the odds and place terms applicable at the time of acceptance. Should a wrong odds or place terms be given in error we reserve the right to settle the bet at the correct odds/place terms that were available at the time the bet was struck.</li>
            </ol>
            <h4>Each-Way Betting</h4>
            <ol>
                <li class="help-li">All bets are settled to win unless 'Each-Way' is selected;</li>
                <li class="help-li">An Each-Way bet is made up of two bets. It contains one bet for your horse to "Win" and a second bet for your horse to be "Placed". Each bet is placed at the stake amount you have entered, so the total cost of an each way bet will be double the amount you entered stake as you are placing two bets;</li>
                <li class="help-li">
                    The "Place" terms will be as advertised for the event. In general, for UK horse racing the 'Place' part of Each-Way bets will be settled using the following 'Place' terms:
                    <ol>
                        <li class="help-li">Less than 5 runners - the place money is invested to win;</li>
                        <li class="help-li">Races of 5, 6 or 7 runners - one 1/4 the odds - first two places;</li>
                        <li class="help-li">All other races of 8 or more runners 1/5 the odds - first three places</li>
                        <li class="help-li">Handicap races with 12 - 15 runners one 1/4 the odds - first three places</li>
                        <li class="help-li">Handicap races with 16 or more runners 1/4 the odds - first four places</li>
                        <li class="help-li">In all races the number of runners will be the number of runners coming                        under starters orders. Bets won't be accepted where the place stake exceeds                        the win stake.</li>
                    </ol>
                </li>
            </ol>
        </li>
    </ol>

    <h3 class="content-item" id="20">
        <strong>Gaelisk spor</strong>
    </h3>
    <ol class="ord-list">
        <li>Outright/Winner insats: Tippa vilket lag som kommer att vinna tävlingen.</li>
        <li>Alla matcher är baserade på ordinarie tid (inklusive övertid). Övertid räknas inte såvida inte specificerat. </li>
        <li>Om något av lagen inte spelar är insatserna ogiltiga. </li>
        <li>Om spelet avslutas före ordinarie tid är insatserna ogiltiga. </li>
        <li>En match som flyttas till en annan dag kommer att vara ogiltig.</li>
        <li>Om en matcharena ändras kommer redan placerade insatser gälla förutsatt att hemmalaget fortfarande är angivet. Om hemma- och bortalaget för en registrerad match ändras kommer insatser placerade på  den ursprungliga registreringen att vara ogiltiga.</li>
        <li>Insatser kommer uteslutande att avgöras på officiella GAA (Gaelic Athletics Association) resultat.</li>
    </ol>
    <h3 class="content-item" id="21">
        <strong>Vintersport</strong>
    </h3>
    <ol class="ord-list">
        <li>
            Outright/Winner insats: Tippa vilket lag som kommer att vinna tävlingen.<li>Alla matcher är baserade på ordinarie tid (inklusive övertid). Övertid räknas inte såvida inte specificerat. </li>
            <li>Om något av lagen inte spelar är insatserna ogiltiga. </li>
            <li>Om spelet avslutas före ordinarie tid är insatserna ogiltiga. </li>
            <li>En match som flyttas till en annan dag kommer att vara ogiltig.</li>
            <li>Om en matcharena ändras kommer redan placerade insatser gälla förutsatt att hemmalaget fortfarande är angivet. Om hemma- och bortalaget för en registrerad match ändras kommer insatser placerade på  den ursprungliga registreringen att vara ogiltiga.</li>
            <li>Insatser kommer uteslutande att avgöras på officiella GAA (Gaelic Athletics Association) resultat.</li>
        </ol>
    <h3 class="content-item" id="22">
        <strong>Vintersport</strong>
    </h3>
    <ol class="ord-list">
        <li>Outright/Winner: Tippa vilket lag/deltagare som kommer att vinna tävlingen. Insatser på deltagare som inte starta kommer inte att betalas tillbaka. </li>
        <li>Vinterolympiad: Tävlingar är officiella efter den ursprungliga medaljceremonin. Eventuella senare ändringar av dessa resultat räknas inte.</li>
    </ol>
    <h3 class="content-item" id="23">
        <strong>Virtual Sports</strong>
    </h3>
    <ol class="ord-list">
        <li>
            <h4>Game Play Rules</h4>
            <ol>
                <li class="help-li">A virtual betting event takes place every 5 minutes.</li>
                <li class="help-li">Bets on the next event are accepted until the "bets closed" message appears on the screen, after which the bet will be allocated to the successive event.</li>
                <li class="help-li">When the event is not specified by the customer, bets are registered on the next event.</li>
                <li class="help-li">Winnings can be collected once the result of an event is displayed on the results screen.</li>
                <li class="help-li">The minimum stake per bet is 50c with a maximum payout for any one customer on any one day of €50,000</li>
                <li class="help-li">A customer who places any bet on these events takes sole responsibility for his actions in placing a bet, and for checking his ticket to ensure it is correctly reflects his chosen bet, and will not 		hold the operator liable in for any loss or damage suffered. The operator will also not be liable for any system malfunction that may result in the nullification, cancellation or refund of a bet at any time.</li>
                <li class="help-li">No horses or greyhounds are scratched from virtual races.</li>
                <li class="help-li">There are no dead heats (position draws) in virtual races.</li>
                <li class="help-li">If any events are cancelled for whatever reason, outstanding bets on the affected events will be paid at settled at 1:1.</li>
                <li class="help-li">Bet types offered may be altered from time to time.</li>
            </ol>
            <h4>Race Event Bet Types &ndash; Single Selection</h4>
            <ol>
                <li class="help-li">
                    <b>Win</b> - Select a runner to finish 1st.
                </li>
                <li class="help-li">
                    <b>Place</b> - Select a runner to finish in 1st, 2nd or 3rd place in a race with 8 runners or more, and 1st, or 2nd in a 6 runner greyhound race.
                </li>
                <li class="help-li">
                    <b>Each-way (“Fractional Place” bet in some fractional odds markets)</b>Select a runner to win or place. This bet consists of two bets on one selection in one event, with the first bet on the runner to 	               			win and the second bet on the runner to place. The place bet pays at a fraction of the win odds as specified on the event data.
                </li>
                <li class="help-li">
                    The Each-Way bet is not offered in most countries. The game system can be configured to set the “place” odds at a fixed proportion of the win odds of the selection as follows:
                    <ol>
                        <li class="help-li">Greyhounds pays 1/5th of win odds.</li>
                        <li class="help-li">Horses pays 1/5th of win odds.</li>
                    </ol>
                </li>
            </ol>
            <h4>Race Event Bet Types - Multiple Selection Combination Odds</h4>
            <ol>
                <li class="help-li">These bet markets carry different terms in different geographical regions. Our data service uses fixed odds (“bookie”) terminology. The system can be configured to display pari-mutuel (“tote”)              terminology on the screen systems and video renders when required. These alternative bet names are shown in parentheses below </li>
                <li class="help-li">
                    <b>Forecast (Exacta)</b> - Select 2 runners to finish 1st and 2nd IN ORDER specified.
                </li>
                <li class="help-li">
                    <b>Combination Exacta</b> - Some bet systems offer a player the option of selecting 2 or more selections to bet that every possible combination of two of the selections may finish 1st and 2nd in               order. So for example; on 2 selections there are 2 bets (1-2, 2-1); on 3 selections there are 6 bets (1-2, 1-3, 2-1, 2-3, 3-1, 3-2); on 4 selections there are 12 bets, on 5 selections there are 20 bets and on 6               selections there are 30 bets etc. This is a bet acceptance system bet that uses the Forecast odds in the feed service. The bet acceptance system works out all combinations.
                </li>
                <li class="help-li">
                    <b>Reverse Forecast (Quinella)</b> - Select 2 runners to finish 1st and 2nd in ANY ORDER.
                </li>
                <li class="help-li">
                    <b>Tricast or Trifecta</b> - Select 3 runners to finish 1st, 2nd and 3rd IN ORDER specified.
                </li>
                <li class="help-li">
                    <b>Combination Trifecta</b> - Some bet systems offer a player the option of selecting 3 or more selections to bet that every possible combination of three of the selections may finish 1st, 2nd and 3rd              in order in an event. So for example; on 3 selections there are 6 bets (1-2-3, 1-3-2, 2-1-3, 2-3-1, 3-1-2, 3-2-1); on 4 selections there are 24 bets; on 5 selections there are 60 bets and on 6 selections there are 120               bets. This is a bet acceptance system bet that uses the Tricast odds. The bet acceptance system works out all combinations.
                </li>
                <li class="help-li">
                    <b>Reverse Tricast or Trio</b> - Select 3 runners to finish 1st, 2nd and 3rd in ANY ORDER.
                </li>
            </ol>
        </li>
    </ol>
    <p style="text-align: right">
        <button type="button" onclick="window.print(); return false" class="button">
            <span class="button_Right">
                <span class="button_Left">
                    <span class="button_Center">
                        <span>Print</span>
                    </span>
                </span>
            </span>
        </button>
    </p>
</div>
