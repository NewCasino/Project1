Transaktionsgräns