﻿<p class="Copy">
			<span class="Hideable">Alla rättigheter förbehålls </span>&copy; 2011&ndash;2012 <a href="/">[metadata:value(/Metadata/Settings.Operator_DisplayNameShort)] Mobile</a>.
		</p>
		<p class="LessEmphasis">
			Oddstjänster som används av  <a href="/AboutUs">[metadata:value(/Metadata/Settings.Operator_DisplayNameShort)] Mobile</a>  tillhandahålls av <a href="http://www.everymatrix.com/">EveryMatrix Ltd</a>. EveryMatrix Ltd. har en klass 2 licens (Nummer LGA/Cl2/497/2008) utfärdad 03.02.2009 av Lotteries and Gaming Authority, Malta, och omfattas av reglering som gäller denna myndighet. Läs mer i <a href="/ResponsibleGaming">Ansvarsfullt spel</a> and our <a href="/TermsConditions">Regler och Villkor </a>.
		</p>

