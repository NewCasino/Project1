Kreditering misslyckades