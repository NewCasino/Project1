﻿ditt bankkonto
