Namn - förnamn