﻿Ditt bankkonto

