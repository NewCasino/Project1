Ogiltig skrill e-postadress.