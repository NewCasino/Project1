Ett konto med samma uppgifter har redan registrerats.