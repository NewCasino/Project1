﻿/game/gamerules.jsp?game=horus&lang=sv