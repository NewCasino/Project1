<p>Hi $FIRSTNAME$,</p><p>Din insättning har blivit nekad. </p><p>Kontrollera den information du matar in och försök igen senare.</p><p>Om du har några frågor tveka inte att kontakta  <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Vänligen,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>