﻿Gå till: 
