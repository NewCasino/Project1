﻿Vänligen fyll i ett giltigt datum
