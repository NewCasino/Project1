﻿Double Exposure Blackjack Serier
