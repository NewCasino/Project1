Uttag av pengar direkt till ditt iDeal-konto