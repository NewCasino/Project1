Erbjudanden