Giltig fr.o.m.