Tillbaka