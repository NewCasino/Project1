﻿Din stad här
