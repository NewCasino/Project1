Mina favoriter