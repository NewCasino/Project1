Formatet i det här fältet är ogiltigt.