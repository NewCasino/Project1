Skicka dina pengar från ditt kreditkort direkt till dina vänner, familj eller företags bankkonton. Det går fort , är enkelt att använda och helt säkert. <br />Vänligen notera att summan som kommer dras förs över i EUR. <br /> Din bank kan komma att ta en växlingsavgift på grund av detta. 