Vänligen infoga sekretesspolicy här[MetaData->PrivacyPolicy].