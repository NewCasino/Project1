﻿ING Bank
