Vänligen välj kompis för överföring