Du har login med fel kontoinformation för många gånger och ditt konto är nu blockad. Vänligen kontakta supporten