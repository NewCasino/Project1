Uttag av pengar direkt till ditt MONETA-konto