﻿Adressrad 2
