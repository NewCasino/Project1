Se till att du noterar dina ändringsuppgifter eftersom du inte kan återgå till den här sidan.