﻿Inloggad
