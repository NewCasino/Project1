Minimalt antal poäng för ansökan: