En 6 månaders själavstängning