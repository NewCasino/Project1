﻿XPro spelande
