﻿Din adress här
