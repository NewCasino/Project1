E-mail addressen kan inte vara tom