﻿Lösenord
