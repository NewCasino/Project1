Se <span class="AlternatesNumber">{0}</span> varianter