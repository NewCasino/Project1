Villkor och bestämmelser