﻿Gör en överföring såsom informationen visas nedanför

