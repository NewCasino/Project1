 värde