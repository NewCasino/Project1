Min favoritfärg?