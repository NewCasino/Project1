﻿/game/gamerules.jsp?game=shvideopokerdw&lang=sv