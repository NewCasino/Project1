﻿Bankkonto valuta
