Uttag av pengar direkt till ditt EPS-konto