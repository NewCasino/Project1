﻿Välj bankkonto