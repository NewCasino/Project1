﻿Ingen tillgänglig bank

