Avgift