﻿Bank 
