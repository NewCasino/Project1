﻿Spela Spel
