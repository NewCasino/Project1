﻿Checkkod
