﻿Maxantal procent
