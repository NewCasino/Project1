﻿Valideringskod
