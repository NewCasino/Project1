Adressen måste bestå av minst 2 tecken