﻿Ta ut direkt till ditt bankkonto
