﻿Min Balansen
