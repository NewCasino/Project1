Betalkort