Betala med textmeddelande