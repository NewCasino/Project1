﻿Your Ukash card