Överför