Starttid