﻿Maxlängd för adressfältet överskriden
