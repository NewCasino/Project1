﻿'marginalBotten'