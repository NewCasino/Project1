Uttag av pengar direkt till ditt AGMO-konto