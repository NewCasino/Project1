Ditt användarnamn innehåller ogiltiga tecken