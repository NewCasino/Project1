﻿Odds Lobby



