﻿/game/gamerules.jsp?game=diamonddogs&lang=sv