﻿<p>Det är inte tillåtet för personer under 18 år att öppna ett konto eller spela på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]. Utöver våra rutiner för slumpmässiga ålderskontroller kommer vi genomföra ålderskontroller på alla kunder vars betalningssätt är tillgängliga för personer under 18 år. Företaget förbehåller sig rätten att begära in dokument som verifierar din ålder, ditt konto kommer att spärras till dess att din ålder har bekräftats.</p>
<p>&nbsp;</p>
<p>Om du delar dator med dina vänner eller familjemedlemmar som är underåriga och du är orolig, överväg en lösning via föräldrakontroll, som är programvaror som ger föräldrar möjlighet att reglera åtkomsten på internet och hindra barns åtkomst till spelsidor.</p>
<p>&nbsp;</p>
<p>Net Nanny&trade; www.netnanny.com</p>
<p>CyberPatrol www.cyberpatrol.com</p>