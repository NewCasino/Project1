﻿Kommande garanteringar
