﻿Slutdatum du har valt är före startdatum
