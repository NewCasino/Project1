﻿Överför pengar med {0}
