﻿/game/gamerules.jsp?game=luckydouble&lang=sv