﻿Vänligen ange ditt namn på kontot
