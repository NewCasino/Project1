Toppkampanj