﻿Klicka för mer information
