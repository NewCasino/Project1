Mitt husdjurs namn?