Ditt Svar