TC nummer