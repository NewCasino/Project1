﻿Vänligen ange din voucherkod
