Internt fel