Sök bord...