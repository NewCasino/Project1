Fortsätt