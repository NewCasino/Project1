Från {0} konto