﻿Neteller(Chile)