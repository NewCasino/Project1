Du har gjort för många inloggningsförsök, så ditt konto har blivit blockerat. Vänta 15 minuter och försök sedan igen.