﻿Förnya Saldon
