﻿Vatican City State