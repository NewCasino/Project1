casinopoäng för frekventa spelare