﻿Vänligen skriv in max belopp


