﻿Belopp som du vill ska dras från ditt konto
