﻿Du kan inte göra en öveföring till dig själv
