﻿/game/gamerules.jsp?game=reelsteal&lang=sv