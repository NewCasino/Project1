Canada dollar