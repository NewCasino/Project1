﻿Fyll i check nummer.