﻿Pris pool
