Adressrad 2 (frivillig)