Alla kampanjer