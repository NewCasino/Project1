[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Registrering bekräftad