﻿Jag vill ha en Bonus. 
