Alla svenska banker