﻿/game/gamerules.jsp?game=halloffame&lang=sv