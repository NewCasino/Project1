﻿TC-NUMMER