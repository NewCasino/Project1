﻿<ol>
        
<li> <strong> Var hittar jag vad kampanjer är i erbjudande? </strong>
<p> Du kan se alla aktuella erbjudanden genom att klicka på vår. [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] kampanjer fliken </p>
</li>

<li> <strong> Kan jag spela alla hemsidan spel när jag tar en bonus, eller finns det några begränsningar på vilka spel jag kan spela? </strong>
<p> Vänligen kontrollera villkoren för bonus och om du är osäker kontakt. [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] kundsupport </p>
</li>


<li> <strong> Hur kontrollerar jag att jag har uppfyllt kraven för en befordran? </strong>
<p> Du kan kontrollera dina framsteg genom att klicka på "Mitt konto" och sedan på vänster du klickar på mitt sport-konto, då aktiva kampanjer. </p>
</li>


<li> <strong> Vilka skäl skulle jag vara sjönk för en befordran? </strong>
<p> Några av de kampanjer kommer att vara berättigade endast för personer från vissa länder och vissa kunder som använder specifika betalningsmetoder. Det kan finnas begränsningar för länkade konton och missbruk av [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] kampanjer, för rådgivning, kontakta [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] Kundtjänst på <a href = "mailto: [Metadata: htmlencode (/Metadata/Settings.Email_SupportAddress)]" target = "_blank"> [Metadata: htmlencode (/Metadata/Settings.Email_SupportAddress)] </a> </p>
</li>
  

</ol>

<p style="text-align:right">
     <button type="button" onclick="window.print(); avkastning false" class="button">
         <span class="button_Right">
             <span class="button_Left">
                 <span class="button_Center">
                     <span> Print </span>
                 </span>
             </span>
         </span>
     </knappen>
</p>
