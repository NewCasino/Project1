Ange avsändarens telefonnummer.