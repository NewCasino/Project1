Vinstsatsers