Ange din e-postadress så skickar vi ett e-postmeddelande med anvisningar om hur du återställer ditt lösenord.