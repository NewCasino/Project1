﻿Belopp som du vill överföra till kortet {0}
