﻿Inbetalning med TLNakit
