Din begäran om tillbakarullning av uttag kan inte handläggas för närvarande.