﻿/game/gamerules.jsp?game=lrroulette2adv&lang=sv