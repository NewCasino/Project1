﻿/game/gamerules.jsp?game=deuceswild100&lang=sv