﻿Pågående
