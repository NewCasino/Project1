﻿CEPBank
