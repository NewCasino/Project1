﻿Du har nått maxantal registrerade kort. För mer info besök vår <a href="/Help">hjälpsektion</a>
