Du kommer inte kunna logga in förrän {0}, är du säker på att du vill fortsätta?