﻿Du måste endast ange nummer i clearingnummersfältet. Vänligen försök igen.
