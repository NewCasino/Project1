Uttag direkt till ditt iDeal konto