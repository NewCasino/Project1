﻿Vinst
