Uttag direkt till ditt VISA kort.