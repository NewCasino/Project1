﻿<style type="text/css">
.limit-overlay{display:none; position: fixed; top: 0; left: 0; z-index: 999998; background: #000; background:  rgba(0,0,0,0.8); filter: alpha(opacity=80);}
.limit-wrap{display:block; width:90%; height: auto;color:#fff; background: #222; border:2px solid #999999; position: fixed; top: 100px; left: 5%; z-index: 999999; }
.limit-box{display: block; margin: 30px auto;}
.limit-box h2{display: block; font-size: 24px; font-weight: bold; text-align: center; margin-bottom: 40px;}
.limit_item{display: block; font-size: 16px; line-height: 20px; margin: 12px 0; text-align: left;}
.limit_item label{margin-left: 20px;}
.limit-buttons{display: block; margin: 30px auto 0;text-align: center;}.limit_type{display: none;}button.limit-button.button {padding: 5px 10px;}
 @media only screen and (max-width: 380px){
.limit-wrap{width:95%;margin-left:2%;left: 0%;}}</style>
