Kortnummer