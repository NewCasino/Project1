﻿Lösenordet måste innehålla minst 7 tecken