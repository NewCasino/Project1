<p> Hej $FIRSTNAME$, </p> Detta automatiserade e-post är ett kvitto på din insättning som bearbetades på uppdrag [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] av EveryMatrix Ltd, betalningsoperatören för [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] hemsida, du kommer att se EveryMatrix på ditt kort eller kontoutdrag. Dina transaktioner är enligt nedan </p> <ul> <li> <strong> Transaction ID </strong>:. $TRANSACTION_ID$ </li> <li> <strong> Datum tid </strong>: $TRANSACTION_ID$ </li> <li> <strong> Webbplats </strong>: $TRANSACTION_ID$ </li> <li> <strong> kvitto </strong>:.  En print screen av ditt kvitto har bifogats </li> </ul > <p> om du har någon fråga angående denna insättning, vänligen kontakta <a med angivande av numret transaktions-ID </p> Hälsningar, <br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]. laget </p> <p>$SCREENSHOT$</p>