Den här transaktionen har slutförts.