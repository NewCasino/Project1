Turkiet lira