Du loggar in från ett land som vi inte tillåter. Vi kommer inte kunna slutföra din registrering.