Fel, det här spelet kan inte spelas i riktiga pengar-läget!