﻿Användarinformation
