Kära $USERNAME$, <br /><br />Syftet med detta e-mail är att bekräfta att din period av 30 dagars självutslutning nu har gått ut och alla funktioner är nu tillgängliga. <br /><br />Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Vänliga Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>