Bonusen har inte aktiverats