Tillåt inte mig att logga in under de nästkommande 7 dagarna