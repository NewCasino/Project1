﻿Väntande
