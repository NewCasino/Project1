Hämtar...