mycket populär