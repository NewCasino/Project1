Ansvarsfullt Spelande