﻿Överför till en vän
