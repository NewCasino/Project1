﻿/game/gamerules.jsp?game=beetle&lang=sv