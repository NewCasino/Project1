﻿Köp in
