﻿Första avlöningsgskravet
