Överföring mellan konton