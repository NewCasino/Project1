﻿/game/gamerules.jsp?game=devil&lang=sv