Valideringskod krävs.