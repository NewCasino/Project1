Ändra lösenord