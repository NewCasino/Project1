﻿You are not eligible to use instaCASH. Please do not enter your bank account information.