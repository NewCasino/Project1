Ny flik