﻿Visa spel i listvy