﻿Läs mer om FPP
