﻿Insättning
