Befintligt kort