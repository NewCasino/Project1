﻿VISA (med GPaySafe)


