Förverka