Du har kopplats från eftersom någon har loggat in med ditt konto från en annan plats.

Om det skett utan ditt godkännande, kan någon ha stulit ditt lösenord och vi rekommenderar att du byter ditt lösenord omedelbart.