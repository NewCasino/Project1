﻿Betsoft spelning
