Alla Spel