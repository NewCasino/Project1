Registreringen är nu slutförd.