﻿PAGOFACIL