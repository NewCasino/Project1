﻿Självexkludera i 6 månader
