﻿/game/gamerules.jsp?game=lrscratchticket&lang=sv