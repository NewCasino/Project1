Startat