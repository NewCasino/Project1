﻿/game/gamerules.jsp?game=hrblackjackpntn&lang=sv