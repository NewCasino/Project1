Kroatien kune