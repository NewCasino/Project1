﻿Vänligen ange ditt användar-ID
