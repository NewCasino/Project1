﻿Speltyp
