Kom ihåg 1 månad