Betala via textmeddelande.