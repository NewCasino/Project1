﻿Upprepa ditt lösenord här
