﻿Muut pelit
