﻿Anmäl dig nu!
