<p>Hej $FIRSTNAME$,</p><p>Tack för att du registrerar dig med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], ditt konto ($USERNAME$) har skapats men innan du kan använda det måste du aktivera ditt konto.</p><p>För att aktivera ditt konto, vänligen klicka på länken nedan, om inget händer, kopiera länken och klistra in den i ett nytt fönster.</p><p><a href="$ACTIVELINK$">$ACTIVELINK$</a></p><p>Om du inte registrerat dig med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], vänligen ignorera detta mail eller informera <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p><p>Tack för din registrering hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]!</p><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>