﻿du kan sätta en så kallad Reality Check som dyker upp på din skärm innan du börjar spela och innebär att det kommer att synas hur länge det har gått sedan du har satt igång med att spela.
