﻿Uttag till
