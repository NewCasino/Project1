﻿Jag är inte tillfredställd med hemsidan
