﻿Direkt banköverföring
