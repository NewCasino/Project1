﻿<p>Hej $FIRSTNAME$,</p>
<p>Du har begärt [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] ändring av din e-postadress.</p>
<p>För din egen säkerhet måste du verifiera din nya e-postadress. För att göra det, klicka bara på länken nedan:</p>
<p><a href="$ACTIVELINK$">$ACTIVELINK$</a></p>
<p>Om länken inte fungerar, kopiera och klistra in länken direkt i din webbläsare.</p>
<p>Om du inte har begärt ändring av din e-postadress, bortse från det här e-postmeddelande eller meddela oss på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p>
<p>Vänliga hälsningar, <br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundtjänstteamet</p>