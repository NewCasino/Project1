Du dirigeras om till {0} sidan, för att insättningen ska slutföras