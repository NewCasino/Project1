﻿Sätt insättningsgräns