Direkt e-banker