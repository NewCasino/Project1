﻿<img src="/Views/Shared/_files/Casino/thumbnail_placeholder.png" />
