Ogiltigt födelsedatum.