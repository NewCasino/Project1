Inloggningen misslyckades. Kontrollera ditt användarnamn och lösenord.