﻿Din e-postadress här
