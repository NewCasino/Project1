Ange skrill e-postadressen.