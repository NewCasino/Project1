Fyll i en IPS token, och för över pengar till den nya kupongen.  