Affiliate-avgift