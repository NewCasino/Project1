Uttag av pengar direkt till ditt TELEINGRESO-konto