﻿Konfiskera alla pengar på utgång
