Felaktig moneybookers e-post adress