Tillåt inte mig att logga in under de nästkommande 6 månaderna