Skickar