Ditt förnamn innehåller otillåtna tecken