﻿<p>Hej $FIRSTNAME$,</p>
<p>Tack för att du registrerar dig hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], ditt konto ($USERNAME$) har skapats och du måste aktivera ditt konto innan du kan använda det.</p>
<p>För att aktivera ditt konto, klicka på länken nedan, om den inte fungerar, försök kopiera och klistra in länken i din webbläsare.</p>
<p><a href="$ACTIVELINK$">$ACTIVELINK$</a></p>
<p>Om du inte har registrerat dig hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], bortse från det här e-postmeddelandet eller meddela <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a></p>
<p>Tack för att du registrerar dig hos [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]!</p>
<p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet</p>