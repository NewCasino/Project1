Mån