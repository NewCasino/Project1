﻿No changes detected