Vänligen ange din stad