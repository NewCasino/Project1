﻿Neteller(Slovakien)
