Bonustyp