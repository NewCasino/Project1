Generellt