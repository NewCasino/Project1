﻿Inbetalning
