﻿Vänligen skriv in ditt bankkontonummer.
