Vänligen fyll i Ukash nummer