Du måste logga in för att spela spelet.