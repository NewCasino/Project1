﻿Februari