Avsändarens TC-nummer