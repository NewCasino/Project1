Ja tack, skicka mig e-mail med nyheter och erbjudanden