﻿Neteller(Hungary)