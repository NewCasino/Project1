﻿Maxlängd av beskrivning är 100 ord. 
