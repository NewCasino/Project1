﻿Setup