Det nya lösenordet kan inte vara samma som det gamla.