Betala per telefon (Kanada)