﻿Till din väns konto


