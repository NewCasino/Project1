﻿Din födelsedag här (DD/MM/YYYY)
