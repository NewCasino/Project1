﻿Gå till hemsidan

