De nästkommande 30 dagarna