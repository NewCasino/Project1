Övrigt