﻿/game/gamerules.jsp?game=lrhilo&lang=sv