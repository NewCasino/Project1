﻿Mobilbetalning
