﻿/game/gamerules.jsp?game=piratesgold2&lang=sv