﻿Net Underhållning
