﻿För att debiteras från kortnr..{0}