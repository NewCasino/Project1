﻿Lägg [metadata:value(/Metadata/Settings.Operator_DisplayName)]till startskärmen!
