Ange captcha.