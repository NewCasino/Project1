Ditt svar måste innehålla minst 2 tecken