﻿Cool-off för 30 dagar
