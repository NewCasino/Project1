Jag vill inte ha någon bonus