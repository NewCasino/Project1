﻿/game/gamerules.jsp?game=lrblackjackdblex&lang=sv