Voucher-numret består av 16 siffror.