﻿HiLo Switch Serier
