﻿Clearingsnummer

