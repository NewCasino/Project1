﻿Odds
