﻿Från {0}