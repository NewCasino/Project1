﻿/game/gamerules.jsp?game=hrblackjackmini&lang=sv