spela på skoj