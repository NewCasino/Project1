﻿/game/gamerules.jsp?game=jacksorbetter1&lang=sv