(uttag endast via banköverföring)