augusti