Vinnare just nu!