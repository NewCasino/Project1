Slutför den här transaktionen i det nya fönstret som öppnats.