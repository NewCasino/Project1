﻿Transaktionshistorik
