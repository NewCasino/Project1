﻿Ogiltig CPR


