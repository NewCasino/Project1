﻿Filtrera