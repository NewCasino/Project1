﻿Slutdatum