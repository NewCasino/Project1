Sidkarta