Användarnamnet är redan taget, välj ett annat