Uttag av pengar direkt till ditt Trustly-konto