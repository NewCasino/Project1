﻿<ol>
        
<li> <strong> Var är din webbplats baserad? </strong>
<p> Vår webbplats är baserad på Malta. </p> </li>

<li> <strong> Är din webbplats licensierat? </strong>
<p> Ja vi har ett giltigt EU-licens för sportsbetting, casino och poker. </p> </li>

<li> <strong> Hur säker är min kreditkortsinformation? </strong>
<p> [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] använder de mest avancerade data krypteringsteknik för att garantera att din information är endast tillgänglig för ett fåtal utvalda inom [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] familj. Vi krypterar all din information med hjälp av internationellt accepterade industristandarder SSL krypteringsalgoritmer. Det innebär all information går fram och tillbaka,. Från din adress, till de kort du håller behandlas är skyddad med samma mått av trygghet en bank skulle använda </p> </li>

<li> <strong> Hur vet jag min ekonomiska information är säker? </strong>
<p> [Metadata: htmlencode (/Metadata/Settings.Operator_DisplayName)] krypterar all din information med hjälp av internationellt accepterade industristandarder SSL krypteringsalgoritmer. Det innebär all information går fram och tillbaka,. Från din adress, till de kort du håller behandlas är skyddad med samma mått av trygghet en bank skulle använda </p> </li>

<li> <strong> Hur vet jag mina pengar är säkra? </strong>
p Alla klientmedel hålls i en separat klient förtroende konto Bank of Valletta. Detta är i överensstämmelse med lotterilagen och förordningar Gaming Malta med vilka vi är licensierade. Klientmedel är helt "öronmärkta" från företagets medel och hålls säkert på detta sätt för att säkerställa att kundernas medel hålls tryggt och finns alltid tillgängliga för klienter. </P> </li>

</ol>
