﻿Ange belopp här
