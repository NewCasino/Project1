﻿Senaste betalkort
