Ett fel inträffade.