﻿Pontoon Serier
