AGMO är ledare inom regional online betalning i CEE regionen. 