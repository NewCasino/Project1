Inga meddelanden 