Ditt efternamn innehåller ogiltiga tecken