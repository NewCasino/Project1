Visa alla tillgängliga spel