﻿                <span class="BannerImg">&nbsp;</span>
                <div class="BannerText">
                    <strong class="MainBannerText">Exclusive Turkish Blackjack tables every day from 8 to 10 pm UCT</strong>
                    <span class="SecondBannerText">Class aptent taciti sociosqu ad litora torquent per conubia nostra, per inceptos himenaeos. Donec malesuada vitae purus non sollicitudin. Phasellus orci augue, porttitor at nunc a, tempor molestie arcu. Quisque ac diam eget neque aliquam consequat at non nunc. </span>
                </div>
