﻿Lägsta insättningsbelopp
