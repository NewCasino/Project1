﻿Jacks or Better -sarja
