﻿Transaktion från spelare {0}