﻿TILLGÄNGLIGA BONUSAR