﻿Endast nummer och / är tillåtet. Vänligen använd punkt för decimaltecken och fyll i nummer utan formatering.
