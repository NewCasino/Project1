﻿Adress linje 2
