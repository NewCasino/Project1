﻿Bonus Bidrag
