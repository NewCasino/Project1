Kampanjlista