Sportbonus Villkor och bestämmelser