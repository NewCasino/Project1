Mottagarens turkiska ID-nummer