﻿Inloggningen misslyckades. Du har valt att självexkludera dig från spelandet till {0}, var god och kontakta kundtjänst efter detta datum.
