valda