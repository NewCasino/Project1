﻿/game/gamerules.jsp?game=allamerican1&lang=sv