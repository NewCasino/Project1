﻿Plånbok
