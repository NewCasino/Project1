﻿Insättning med <span>{0}</span>
