﻿Neteller(Turkiet)
