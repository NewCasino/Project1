Sortera