﻿Överför från ditt {0} konto
