Uttaget kommer processas så fort som möjligt