Välj en kompis.