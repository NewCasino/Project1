﻿Dubbel Jackpot Poker
