﻿Ta ut direkt till ditt AstroPayCard konto
