﻿Neteller(Sverige)
