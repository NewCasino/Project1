Ukash (av Dotpay)