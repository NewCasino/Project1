﻿Fyll i betalare