Personuppgifter