﻿Formatet i fältet är ogiltigt . ( e.g. AABAFI22 eller NDEAFIHH030 )
