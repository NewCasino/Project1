﻿Van Lanschot
