﻿<p>Hi $FIRSTNAME$,</p>
<p>Din insättning har slutförts</p>
<p>
  <span style="font-size: medium;">
    <strong style="color: #ff3366;">Klicka på "Uppdatera" knappen(NOT the web browser refresh button) överst på sidan för att uppdatera ditt saldo</strong>
  </span>
</p>
<p>
 Om du har några frågor tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.
</p>
<p>
  Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team
</p>


