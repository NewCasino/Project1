﻿<p>Dear&#160; $USERNAME$,<br />
<br />
Du får det här mailet eftersom dina kumulativa uttag har nått 2300 €. Vi är skyldiga att bekräfta din identitet när de kumulativa uttagen har nått 2300€ för att följa maltesiska och europeiska lagar, föreskrifter och riktlinjer för att förebygga penningtvätt och finansiering av terrorism. Alla transaktioner som görs av spelare kontrolleras för att förhindra penningtvätt och all annan olaglig verksamhet. Genom att acceptera Regler & Vilkor tillåter du oss att utföra verifieringar.
<br />
Vänligen skicka legitimation såsom pass eller nationellt ID till <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>. När verifieringen är slutförd, kommer ditt uttag behandlas omedelbart.
<br />Om du inte kan ge dessa bevis, kommer ditt konto bli tillfälligt eller permanent stängt.
<br />
Hälsningar,<br />
[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team
