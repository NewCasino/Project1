﻿Spela på riktigt
