﻿Variabel