Utfärda en IPS-token