Mitt husdjursnamn?