Beskrivning