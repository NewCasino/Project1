﻿Max Belopp


