﻿Välj konto