﻿Tillbaka

