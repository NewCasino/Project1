﻿Öppna visning av spel från {0}