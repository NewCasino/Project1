﻿/game/gamerules.jsp?game=hrblackjackdblex&lang=sv