Registrera ett konto