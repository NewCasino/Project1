﻿/game/gamerules.jsp?game=marbles&lang=sv