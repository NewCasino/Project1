﻿Cool-off för 7 dagar
