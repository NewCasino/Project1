Verifieringskod