﻿/game/gamerules.jsp?game=jokerwild5&lang=sv