[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Live Kasino