﻿Bekräfta lösenord
