Du måste logga in för att ändra din e-postadress.