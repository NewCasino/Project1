i turneringar