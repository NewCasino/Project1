Avbryt Uttag