﻿Emailadress
