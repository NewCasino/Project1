AnvändarID