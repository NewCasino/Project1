﻿Jacks or Better Serier
