﻿Vänligen ange verifieringskoden

