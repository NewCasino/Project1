Befintligt konto