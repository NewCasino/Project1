Denna alias används redan.