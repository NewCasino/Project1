Ange insättningsgräns