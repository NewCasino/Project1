Vänligen ange ditt förnamn