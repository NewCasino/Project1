﻿Fel. Kontrollera dina uppgifter och prova igen
