﻿Välj Debetkonto


