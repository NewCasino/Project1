Slutför