﻿Maxlängd för ortfältet överskriden
