Din nya e-postadress har verifierats och aktiverats.