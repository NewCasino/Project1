﻿Casinospel - FPP-satser