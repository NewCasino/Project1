﻿Bordet är för närvarande stängt. Vänligen återkom mellan {0}. 

