﻿Vänligen välj ett insättningskonto