﻿Öppetider:

