Störst vinnare: