Visa spel med ikoner i ett rutnät