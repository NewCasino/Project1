Verifiera din överföring