﻿Spelkupong
