[Metadata:value(/Metadata/Settings.Operator_DisplayName)], ansvarsfullt spelande