﻿Landfältet får inte lämnas tomt
