Ange börs.