﻿Välj en vän
