Omedelbar