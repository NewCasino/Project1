﻿Självexkludera i 5 år
