﻿Kampanjer - $CATEGORY$
