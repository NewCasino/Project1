Sortera efter populäritet