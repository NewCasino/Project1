﻿Ditt användarnamn här
