Alla jackpottar