﻿SNS Regio Bank
