﻿Konto-ID