Inkorrekt mobilnummer