Ämne