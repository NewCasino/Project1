Alla spel