belopp här