Tillgänglig bonus