Ange TC-NUMRET.