<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Din personliga tidsbegränsning är bestämd till $NYPERIODGRÄNS$ minuter. <br /><br /> Du kan minska din tidsbegränsningomedelbart genom att använda samma meny inom området Ansvarsfullt Spelande på sidan <br /><br /> Om du önskar öka din gräns kommer det ta 7 dagar innan den nya gränsen aktiveras. Perioden om 7 dagar ges för att tillåta dig dig att under tiden ompröva ändringen om så nödvändigt.<br /><br />Vänligen tveka inte att kontakta oss om du har några frågor på<a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet   </p>