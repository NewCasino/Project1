Transaktion ID