﻿Kontakinformation
