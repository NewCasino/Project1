﻿Det gick inte att läsa in balansen, försök igen senare.
