﻿Du behöver logga in för att se din profil