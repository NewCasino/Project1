[Metadata:value(/Metadata/Settings.Operator_DisplayName)] - Ditt konto är blockerat