﻿Hitta en vän genom användarnamnet
