Vinnande spel: {0}