﻿Din väns konto är inaktivt
