Integritetspolicy