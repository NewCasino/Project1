﻿Uttag direkt till ditt UIPAS-konto
