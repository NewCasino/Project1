﻿<img src="//cdn.everymatrix.com/Shared/_files/Deposit/CardGuide_CVCNumber.png" />
<br />
<span>Den består av 3 siffror och finns på baksidan av ditt kort.</span>