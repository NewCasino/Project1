Uttag direkt till ditt EUTELLER konto