﻿Neteller(Frankrike)
