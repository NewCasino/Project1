Vänligen fyll i moneybookers e-post adress