﻿Dölj Vågar
