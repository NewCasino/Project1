﻿[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Din e-postadress har ändrats.