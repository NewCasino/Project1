﻿Transaktionen kunde inte utföras för tillfället
