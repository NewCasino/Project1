Bakåt