Uttag av pengar direkt till ditt TLNakit-konto.