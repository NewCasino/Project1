﻿Steg 1 / 2. Det tar bara två minuter
