TILLGÄNGLIGA BONUS