TransaktionsID