Konto information