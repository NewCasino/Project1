﻿Jag vill inte sätta en gräns just nu
