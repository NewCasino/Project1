Meddelande