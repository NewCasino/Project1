Gräns för sessionstid