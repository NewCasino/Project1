Personligt ID nummer