﻿Användarnamnet måste innehålla minst 4 tecken
