﻿Du måste logga in för att avbryta uttag
