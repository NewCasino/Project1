Att ta från {0}