﻿Ta ut direkt till ditt VISA-kort
