E- {0} postadressen har redan registrerats på {1}, om du vill associera ditt {2} konto med ditt existerande {1} konto ska du logga in här.