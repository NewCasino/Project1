﻿Neteller konto-ID eller E-postadress