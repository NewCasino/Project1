﻿poytapelit

