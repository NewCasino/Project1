﻿Maxlängden för fältet som är avsedd för ditt förnamn är överskriden
