Du kommer inte kunna logga in på ditt vadslagningskonto under avkylningsperioden av 1 år