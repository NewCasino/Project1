ogiltige-mail format