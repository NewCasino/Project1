Meddelandet har skcikats, vi ger dig en återkoppling så snart som möjligt