Uttag av pengar direkt till ditt BOLETO-konto