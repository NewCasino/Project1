Aktivera ditt konto