Om kontanta vinster