﻿Tens eller Bättre Serier
