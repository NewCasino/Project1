﻿Ingen information
