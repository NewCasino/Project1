﻿Mina Spel
