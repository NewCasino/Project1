﻿Ditt lösenord här
