﻿Ta ut dina pengar
