﻿Videopokerit
