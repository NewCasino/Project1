Detta fält är nödvändigt