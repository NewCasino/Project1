Du måste logga in för att kunna spela spelet i riktiga pengar-läge.