﻿Har du inget konto än?
