Se alla kampanjer nu!