﻿Att dras från ditt konto:
