Må