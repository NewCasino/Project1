Prispool