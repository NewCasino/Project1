[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Kontakta oss