﻿/game/gamerules.jsp?game=boombrothers&lang=sv