Vi har även möjlighet att stänga ditt konto permanent: