﻿/game/gamerules.jsp?game=deuceswild1&lang=sv