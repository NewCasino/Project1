Ange ditt förnamn