Ingen sortering av spelen