Lösenordet får inte vara detsamma som användarnamnet.