Utgångsdatum