﻿Vänligen ange din mobil.
