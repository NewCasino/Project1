﻿Skapa konto nu!


