﻿/game/gamerules.jsp?game=jacksorbetter100&lang=sv