Spela LIVE BlackJack nu!