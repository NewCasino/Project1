﻿BankLink (U|NET)