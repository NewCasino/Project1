﻿Bonuserbjudande
