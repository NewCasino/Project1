Betala per telefon (Belgien)