[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Anmälan av ändrad e-mailadress