Vänligen ange valuta