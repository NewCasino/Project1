﻿Har du glömt ditt Lösenord?


