Ikonerna betyder: