﻿Du har blivit frånkopplad för att någon har loggat in med ditt konto från en annan enhet.

Observera om detta inte är medvetet kan någon ha stulit ditt lösenord, vi rekommenderar dig att byta lösenord snarast.

