﻿Trustly (med MoneyMatrix)
