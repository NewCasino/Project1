﻿Casinospel
