﻿[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] - Verifiering av ändrad e-postadress