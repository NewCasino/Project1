Du kan för närvarande inte ändra din e-postadress eftersom ditt konto är inaktiverat. Ett aktiveringsmeddelande har skickats till e-postadressen som du angav vid registreringen. Klicka på länken i aktiveringsmeddelandet för att aktivera ditt konto. Om du inte får aktiveringsmeddelandet, kontakta <a href="mailto:[Metadata:value(/Metadata/Settings.Email_SupportAddress)]">[Metadata:value(/Metadata/Settings.Email_SupportAddress)]</a>.