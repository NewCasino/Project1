﻿CA$ (CAD)
