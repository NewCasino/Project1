Insättning {0} {1} för {2} {3} Bonus