﻿Logga in


