﻿/game/gamerules.jsp?game=voodoo&lang=sv