﻿SWIFT är fel. Du får inte använda det angivna SWIFT-numret.
