﻿Blackjack Progressive US