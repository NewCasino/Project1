﻿Vänligen ange medborgar ID
