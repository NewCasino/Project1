Du kan inte besöka den här sidan på grund av ofullständig profil. Du dirigeras vidare om 5 sekunder, komplettera din profil och försök igen.