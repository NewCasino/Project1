Banköverföring