Konto ID