﻿Klicka <a href="https://www.uipas.com/home/register" target="_blank">här</a> registrera ditt UIPAS konto idag för insättning.
