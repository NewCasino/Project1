﻿Fel
