﻿NEJ
