<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Din personliga förlustgräns är bestämt till $NEWLIMITAMOUNT$ $NEWLIMITPERIOD$. <br /><br /> Du kan minska din förlustgräns omgående genom att använda samma meny på området Ansvarsfullt spelande på sidan. <br /><br /> Om du skulle vilja öka din gräns så tar det 7 dagar innan den nya gränsen aktiveras. 7-dagars perioden ges så att du hart id att tänka över ändringen om så är nödvändigt.<br /><br /> Vänligen tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet Team   </p>