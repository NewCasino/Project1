﻿Hilo Switch Serier
