﻿Valutafältet får inte lämnas tomt
