ange check-numret.