Metoden att betala per telefon är exakt vad det låter som: betala per telefon, och det är också ettlämpligt betalningsätt från en mobiltelefon. Kunderna ringer ett nummer och betalar per minut, eller per samtal. Denna metod av betalning är idealisk för så kallade ”microbetalningar”, och erbjuder en metod av betalning för målgrupper som inte har ett kreditkort eller ett eget bankkonto.