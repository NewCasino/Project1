﻿Domain status was not changed