﻿/game/gamerules.jsp?game=jokerwild50&lang=sv