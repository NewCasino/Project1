﻿Spel
