(Frivillig)