﻿<img src="//cdn.everymatrix.com/_casino/5/5767E9DF8FE4B02067D0419AD4F14BA7.jpg" />
