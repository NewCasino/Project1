﻿(valfritt)
