maj