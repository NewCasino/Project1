﻿Ditt lösenord ska bestå av minst 6 tecken
