Bank transfer