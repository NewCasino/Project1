Du måste logga in för att göra en självuteslutning.