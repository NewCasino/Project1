Klicka på Slutför häri för att uppdatera dina transaktionsuppgifter.