Börs