Riktiga pengar