﻿Nedtrappning under 24 timmar
