Kom inte ihåg