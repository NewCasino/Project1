﻿Du måste ange nummer i kontonummersfältet. Vänligen försök igen.
