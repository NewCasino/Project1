Bonusvillkor och -bestämmelser