﻿
  <h1><a href="/">SMSCoins - zamień SMSa na żetony<span></span></a></h1>
  <div id="content">
    <div class="box" id="zeton5">
      <h2>25 żetonów<span></span></h2>
      <div class="box-content">
        <p class="firstp">Aby otrzymać 25 żetonów o wartości 2,50 zł,</p>
        <p>wyślij sms-a o treści <strong>AP.ZETON5</strong> na numer <strong>75068</strong>. <span>Koszt przesłania wiadomości wynosi 6,15&nbsp;zł brutto.</span> </p>
      </div>
    </div>
    <div class="box" id="zeton6">
      <h2>30 żetonów<span></span></h2>
      <div class="box-content">
        <p class="firstp">Aby otrzymać 30 żetonów  wartości 3,00 zł,</p>
        <p>wyślij sms-a o treści <strong>AP.ZETON6</strong> na numer <strong>76068</strong> <span>Koszt przesłania wiadomości wynosi 7,38&nbsp;zł brutto.</span> </p>
      </div>
    </div>
    <div class="box" id="zeton9">
      <h2>45 żetonów<span></span></h2>
      <div class="box-content">
        <p class="firstp">Aby otrzymać 45 żetonów o wartości 4,50 zł,</p>
        <p>wyślij sms-a o treści <strong>AP.ZETON9</strong> na numer <strong>79068</strong> <span>Koszt przesłania wiadomości wynosi 11,07&nbsp;zł brutto.</span> </p>
      </div>
    </div>
    <div class="box" id="zeton19">
      <h2>95 żetonów<span></span></h2>
      <div class="box-content">
        <p class="firstp">Aby otrzymać 95 żetonów o wartości 9,50 zł,</p>
        <p>wyślij sms-a o treści <strong>AP.ZETON19</strong> na numer <strong>91958</strong> <span>Koszt przesłania wiadomości wynosi 23,37&nbsp;zł brutto.</span> </p>
      </div>
    </div>
    <div class="box" id="zeton25">
      <h2>125 żetonów<span></span></h2>
      <div class="box-content">
        <p class="firstp">Aby otrzymać 125 żetonów wartości 12,50zł,</p>
        <p>wyślij sms-a o treści <strong>AP.ZETON25</strong> na numer <strong>92578</strong> <span>Koszt przesłania wiadomości wynosi 30,75&nbsp;zł brutto.</span> </p>
      </div>
    </div>
  </div>
  <div id="footer">
    <p>Copyrights &copy; 2009 smscoins.net</p>
  </div>
  <p id="footer2"> Usługa działa we wszystkich sieciach polskich operatorów.<br>
    Uwaga! Możesz przesłać jedynie 1 SMS o wartościach 19 i 25 zł w ciągu 20 minut<br>
    oraz 2 SMSy o pozostałych wartościach. </p>
  <p style="text-align:center"> <a href="/">regulamin</a> </p>
