Ogiltigt SWIFT, du kan inte använda vårt exempel-SWIFT.