﻿Singel Blackjack
