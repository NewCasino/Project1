Mitt mellannamn?