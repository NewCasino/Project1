Ämne.