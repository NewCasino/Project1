Laddar...