﻿Withdrawal requires at least one successful deposit