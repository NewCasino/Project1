﻿Vänligen skriv in ett belopp att överföra


