﻿Spelutveckling
