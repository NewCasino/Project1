Sortera spelen efter prioritets- eller alfabetisk ordning.