Din mobil stöds inte av vald bank, du måste uppdatera din mobil för att kunna fortsätta insättningen.