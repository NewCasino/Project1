Du kan inte göra en insättning för att ditt konto är inaktiverad Ett aktiveringsmail har skickats till din e-post då du registrerade kontot.Vänligen klicka på länken i mailet för att akitvera ditt konto. Om du inte har fått aktiverings mailet så kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.