Ange ditt bankkontonummer.