Vänligen fyll i lösenord.