﻿/game/gamerules.jsp?game=hilo2-3c&lang=sv