Procentuellt maxbelopp