﻿Säkerhetskoden krävs
