﻿Markera rutan!
