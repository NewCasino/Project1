Kortinnehavarens namn är obligatorisk.