Uttag av pengar direkt till ditt Maestro-kort.