Mrs