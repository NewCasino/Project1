Direktbank