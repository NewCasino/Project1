Om detta inte stämmer och du kom hit genom att klicka på en länk som vi har skickat till dig, kan länken vara för gammal nu.