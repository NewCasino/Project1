Du kommer inte kunna logga in på ditt vadslagningskonto någonsin igen