Klicka för att visa guiden.