Snabbregistrering med