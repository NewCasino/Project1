﻿Triodos Bank
