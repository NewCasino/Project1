Summa debiterat från ditt {0} konto