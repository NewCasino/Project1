Direktdebitering från ditt bankkonto.