Du måste logga in för att se den här sidan