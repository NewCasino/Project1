Uttag direkt till dittVISA electron kort.