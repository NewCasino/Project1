﻿Your request could not be completed. An unknown error has occurred. Please try again. Email {email address} if you continue to receive this error.