Skicka nu