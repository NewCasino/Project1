﻿//static.gammatrix-dev.net/MobileShared/_files/top-logo@2x.png

