﻿Din mailadress här
