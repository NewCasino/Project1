﻿/game/gamerules.jsp?game=lrbaccarat2&lang=sv