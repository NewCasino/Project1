﻿Du måste vara inloggad för att kunna överföra pengar.
