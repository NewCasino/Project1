Ange ditt lösenord.