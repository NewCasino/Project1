Avsändarens TC nummer