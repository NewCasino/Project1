﻿Cuenta Digital