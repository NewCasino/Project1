﻿Transaction Historia
