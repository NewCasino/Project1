﻿Vänligen fullfölj överföringen i fönstret som öppnas upp
