﻿Augusti