﻿Din väns användarnamn
