﻿Var vänlig och se till att den valda valutan ovan och ”Ukash värde” nedan är i samma valuta och samma mängd som ditt Ukash kort.
