﻿AU$ (AUD)
