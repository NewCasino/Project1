﻿Friesland Bank
