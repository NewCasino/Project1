Ange ditt konto-ID