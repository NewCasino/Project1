Lägg till i Favoriter