Betala per telefon (USA)