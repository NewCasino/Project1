Daglig gräns