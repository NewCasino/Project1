﻿Har du inget NETeller konto? Klicka <a href="/Deposit/NetellerQuickRegister">här</a> för att öppna ett.
