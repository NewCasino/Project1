Mobilsida