﻿Öppna konto
