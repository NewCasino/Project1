﻿Du spelar på skoj. <a class="Button IncentiveButton" href="#" title="Logga in eller öppna ett konto nu!">Spela med riktiga pengar</a>