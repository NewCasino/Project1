Se nästa spelsida