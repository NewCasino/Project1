Belopp som dras från {0} konto.