﻿Ditt svar här
