﻿Utfärdare
