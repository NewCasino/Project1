Namn - Förnamn