﻿Arvonta
