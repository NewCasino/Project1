Språk