﻿Max.allowed attachment number ({0}) exceeded