Välj konto för debitering