Din insättning av pengar lyckades