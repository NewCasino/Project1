﻿Existerande kort
