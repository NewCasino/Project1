﻿Ogiltigt konto ID.
