Debiterad avgift