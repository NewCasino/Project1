﻿All American Series