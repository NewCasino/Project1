﻿Spela för riktiga pengar

