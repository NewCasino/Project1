Markera markeringsrutan!