﻿/game/gamerules.jsp?game=fortuna&lang=sv