﻿Tillåta erbjudanden via SMS
