﻿Vänligen ange ditt efternamn
