Nigeria naira