Annullerad