Ange belopp