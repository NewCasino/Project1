Välj ditt användarnamn