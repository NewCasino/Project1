﻿The account number is invalid