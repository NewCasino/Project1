Mitt konto