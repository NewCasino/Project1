﻿Maj