Ange din skattekod