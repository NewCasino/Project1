﻿Lösenord:


