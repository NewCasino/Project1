Ditt Secure ID måste vara minst 6 tecken