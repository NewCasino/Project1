<p>Kära $USERNAME$,</p><br /> Tack för att du kontaktat [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]<br /><br /> Syftet med detta e-mail är att bekräfta att din personliga tidsbegränsning ($PERIODSGRÄNSER$ minuter) kommer att tas bort på $LIMITEXPIRYDATE$. <br /><br /> Var vänlig, tveka inte att kontakta oss om du har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p><br /> Vänliga hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kundsupport teamet</p>