Vänligen fyll i avsändarens telefonnummer