Uttag av pengar direkt till ditt NEOSURF-konto