Välj ett spel: