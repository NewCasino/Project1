﻿other-games
