Ta bort {0} från dina favoriter