Rum