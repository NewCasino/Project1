﻿Riktig brasilianska