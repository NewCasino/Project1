﻿i-BANQ användar-MID är fel
