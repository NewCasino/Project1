﻿Alternativa betalningsväxel
