Dölj knappen för öppning av slumpmässigt bord