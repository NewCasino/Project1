Min mammas flicknamn?