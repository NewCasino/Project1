﻿/game/gamerules.jsp?game=junglegames&lang=sv