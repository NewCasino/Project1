﻿Jag vill ha en bonus.
