Pågår