﻿Titel måste anges
