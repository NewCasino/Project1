Bonusnamn