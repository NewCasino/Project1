﻿Avgift