﻿Gå tillbaka
