﻿Ditt ämne här
