Max.  {0} {1:N0}