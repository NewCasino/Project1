﻿XPro Spelning
