﻿Användarnamn:
