E-mailadressen är inte tillgänglig eller har redan använts av någon annan, var vänlig prova en annan e-mail.