﻿IGT Spel
