Du måste logga in för att visa din profil.