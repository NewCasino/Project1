﻿Ditt efternamn här
