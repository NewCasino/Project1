Bingo-rum