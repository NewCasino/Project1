﻿Fyll i banknamn