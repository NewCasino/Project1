﻿Sätt din gräns
