Summa