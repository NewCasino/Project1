Du kommer inte att kunna logga in på ditt bettingkonto under uppehållsperioden på 7 dagar