﻿Vi har för närvarande inga aktiva kampanjer för detta avsnitt. Kom tillbaka senare.
