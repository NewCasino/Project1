﻿Meddelande sänt

