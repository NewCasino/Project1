Stad måste innehålla minst 2 tecken