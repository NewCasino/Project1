﻿<p class="ATHP">Tap the <span class="ATHIcon">Lägg till startskärmen</span> ikonen nedan och välj "Lägg till på hemskärmen".</p>
