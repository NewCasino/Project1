﻿Land Blokerat
