﻿Användarnamn
