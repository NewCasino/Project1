﻿Personal ID nummer