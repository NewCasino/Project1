Teoretisk utbetalning