﻿Meny
