Behandlas