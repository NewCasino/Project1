﻿Videopokerit

