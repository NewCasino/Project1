Fel e-postformat.