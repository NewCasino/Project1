Välj lösenord