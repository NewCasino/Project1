﻿Neteller(Japan)