﻿Du har en pågående insättningsförfrågan, var god och vänta tills denna har godkänts av vårt team. För detaljer, kontakta live support.
