Dina gränser