Omedelbart