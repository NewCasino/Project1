﻿Sätt en spelsessionsbegränsning
