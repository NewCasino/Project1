Bankkod/typkod