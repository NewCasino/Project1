Ange bankkoden.