Du måste bekräfta att du är minst {0} år