﻿You have requested an amount below {$}. Please try again.