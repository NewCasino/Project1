Använd senast