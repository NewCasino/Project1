﻿Väntande uttagsförfrågan
