﻿Smart underhållning
