﻿/game/gamerules.jsp?game=deuceswild50&lang=sv