Processen har lyckats!