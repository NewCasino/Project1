Spela {0} på skoj