﻿Observera att din insättning behandlas av EveryMatrix Ltd, betalningshandläggare för [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] webbsida, kommer du att se Internetbetalning på ditt kontoutdrag.