Ange din stad/ort