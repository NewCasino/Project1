Uttag direkt till ditt Trustly konto