Du måste logga in för att ange en insättningsgräns.