Visa spel i listvy