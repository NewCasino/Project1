Vänligen välj din säkerhetsfråga