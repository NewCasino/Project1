Kopiera