﻿OS Spel
