﻿Validation kod är obligatorisk.