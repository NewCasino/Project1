Ange din e-postadress så skickar vi ett e-postmeddelande med ditt användarnamn.