Landet där du bor