Ange mottagarens TC-nummer.