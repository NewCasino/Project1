﻿Pågående