Max summa