Sö