﻿Tillgången till kontot har nekats då du har självexkluderat dig i ROFUS.

