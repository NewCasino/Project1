﻿Konto