Hemlig access-kod