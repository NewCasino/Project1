Vänligen välj ett kort