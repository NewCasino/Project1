﻿/game/gamerules.jsp?game=letitride2&lang=sv