﻿/game/gamerules.jsp?game=allamerican50&lang=sv