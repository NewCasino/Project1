﻿Logga ut
