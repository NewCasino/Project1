﻿Vänligen kontakta support om du har frågor
