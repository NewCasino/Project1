Gör ett uttag direkt till ditt Balotokonto