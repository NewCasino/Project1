﻿Kommande freerolls
