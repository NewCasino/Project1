Laddar…