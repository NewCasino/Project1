﻿nära:stäng detaljer
