﻿/game/gamerules.jsp?game=fiftyhvideopokerdw&lang=sv