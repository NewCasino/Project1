Du kommer aldrig mer att kunna logga in på ditt bettingkonto