﻿Risk Rejection due to IP Country check. For further assistance, please contact service@click2pay.com