﻿
<ol>
<li> <strong> Jag har glömt mitt användarnamn och lösenord , vad gör jag ? </strong >
<p> Ange ett felaktigt lösenord kan ofta resultera i en " inte kan validera lösenord " kod . Eftersom lösenord är skiftlägeskänsliga , kontrollera din Caps Lock är avstängd . Om dina problem kvarstår , välj " glömt lösenord "-knappen och ett nytt lösenord kommer att utfärdas till den e - postadress som anges på [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] . Konto </p >
</li >

<li> <strong> Vem ska jag kontakta om jag har frågor om mitt konto ? </strong >
<p> Vänligen kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] Kundtjänst <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank"> [ Metadata : htmlencode (/Metadata/Settings.Email_SupportAddress ) ] </a > </p >
</li >

<li> <strong> Vad gör jag om jag inte längre vill använda mitt konto ? </strong >
<p> för att stänga kontot maila [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] Kundtjänst på < a href = " mailto : [ Metadata : htmlencode (/Metadata/Settings.Email_SupportAddress ) ] " target = " _blank " > [ Metadata : htmlencode (/Metadata/Settings.Email_SupportAddress ) ] </a > </p >
</li >

<li> <strong> Hur ändrar jag mitt lösenord ? </strong >
<p> Du kan ändra lösenordet med hjälp av den bortglömda - lösenord <a href="/ForgotPassword" target="_blank"> länk </a > på toppen av alla [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] sidor . </p>
</li >

<li> <strong> Hur ändrar jag min registrerade e-postadress ? </strong >
<p> Vid denna tid kan du inte själv ändra din e-postadress , men om du kan visa goda skäl för den e-postadress ändras , vänligen kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] Kundsupport för eventuella ändringar i dina kontouppgifter . Vänligen kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank"> [ Metadata : htmlencode (/Metadata/Settings.Email_SupportAddress ) ] </a > </p >
</li >

<li> <strong> Finns det något sätt jag kan kolla mitt konto aktivitet ? </strong >
<p> Du kan kontrollera ditt konto aktivitet genom att gå till " Mitt konto " när du har loggat in , eller så kan du kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] . Kundtjänst för information </p >
</li >

<li> <strong> Är det möjligt att ändra mitt användarnamn ? </strong >
<p> Du kan inte ändra ditt spelarnamn när du har skickat till din [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] konto . Detta är av säkerhetsskäl sedan ändra spelarens namn kan störa systemet data och höjer säkerhetsvarningar . </P >
</li >

<li> <strong> Vem kan jag kontakta om jag tror att jag har ett problem med mitt spelande ? </strong >
<p> delta i online gaming är spännande , roligt och potentiellt lönsamma för dem som valde att spela . Men [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] är medveten om möjligheten av spel missbruk och de återverkningar det kan ha på en individ . På grund av detta , [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] tar alla försiktighetsåtgärder för att säkerställa att våra produkter och tjänster används endast av dem som har laglig rätt att göra det . Under inga omständigheter är några spelare tillåts att spela för riktiga pengar om de inte uppfyller åldersgräns på 18 eller standarden laglig ålder för att delta i online- spel i det land där de är bosatta . </P >
</li >

<li> <strong> Vad händer efter min tid är upp ? </strong >
<p> När tidsgränsen du valt för egen uteslutning är upp kan du kontakta [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] Kundtjänst för att öppna ditt konto </p > .
</li >

<li> <strong> Hur kan jag själv utesluta ? </strong >
<p> Du kan själv utesluta genom att gå in i din [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] konto , där du kommer att se själv axclusion fliken när du trycker på Block mitt konto knapp , kommer du automatiskt logga ut den [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] webbplats . Den inloggningen kommer då endast att vara möjligt efter utgången av den tillgång preskriptionstiden du valt . </P >
</li >

<li> <strong> Kan jag avboka det ? </strong >
<p> Du kan inte öppna ditt konto förrän den tidsperiod du valt för egen uteslutning är klar . </p >
</li >

<li> <strong> Jag får inte ett svar på mina frågor när jag e - post Support Team ? </strong >
<p> Vi strävar efter att svara på alla kundservice e-post inom 24 timmar . Som en del kräver mer detaljerat och utredningen av en fråga , kan svarstiden variera beroende på vilken typ av din förfrågan . Du kommer att få ett e - post bekräftelse från [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] när vi har mottagit din förfrågan , så att du vet att vi arbetar på ett svar . Om du upptäcker att du inte får den bekräftelse via e - post omedelbart efter att skicka din förfrågan föreslår vi att du har en titt i din skräppostmapp . [ Metadata : htmlencode (/Metadata/Settings.Operator_DisplayName ) ] . Inte engagera sig i handlingen att skicka oönskad e-post men några aggressiva postfilter kan ibland identifiera våra e-postmeddelanden som spam och behandla dem som sådana </p >
</li >
</ol >

<p style="text-align:right">
    <button type="button" onclick="window.print(); avkastning false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span> Print </span >
                </span >
            </span >
        </span >
    </knappen >
</p >

























































 


 
 

 

 


 
 

 

 


 
 

 

 






Google Translate for Business:Translator ToolkitWebsite TranslatorGlobal Market Finder









Turn off instant translationAbout Google TranslateMobilePrivacyHelpSend feedback

