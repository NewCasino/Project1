Välj din valuta