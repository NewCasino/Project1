﻿Andra Spel
