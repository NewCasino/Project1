﻿The requested functionality is not available or not supported in the current configuration.