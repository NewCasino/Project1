Alla medel kommer att förverkas i enlighet med de Villkor och bestämmelser som du har godkänt, är du säker på att du vill fortsätta?