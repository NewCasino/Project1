Länken har utgått eller är ogiltig