Blocka ditt konto