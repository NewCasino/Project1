﻿Ditt bankkonto
