Ekonomi