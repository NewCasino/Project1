﻿Adressinformation
