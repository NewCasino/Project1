﻿Spela i vårt Casino
