Ange ett nytt lösenord