Repetera lösenordet