Bonuskoden har godkänts!