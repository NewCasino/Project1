Största jackpots