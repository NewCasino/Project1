﻿EcoCard