﻿Mitt Saldo...
