I menyn nedan kan du välja hur mycket du vill sätta in på ditt konto per dag, per vecka eller per månad. Dessa gränser är oberoende av gränserna eller de lägsta gränserna som erbjuds via metoderna på insättningssidan. När en gräns har angetts, får du ett bekräftelsemeddelande via e-post. Du kan minska din gräns när som helst via den här menyn. Men, om du vill återställa dina gränser (vilket kan göras med knapparna nederst på sidan) tillämpas en 72-timmars väntetid (den här perioden ger dig tid att fundera över din ändring). Observera att den här insättningsgränsen är baserad på ditt netto.