Du måste logga in för att överföra pengar.