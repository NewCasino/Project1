﻿Registrera
