Stad/ort