﻿/game/gamerules.jsp?game=hrletitride2&lang=sv