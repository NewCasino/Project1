﻿Dubbel Bonus Poker
