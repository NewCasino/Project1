﻿Denna fält är obligatorisk