﻿/game/gamerules.jsp?game=jokerwild10&lang=sv