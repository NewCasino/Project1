﻿Självavstängning