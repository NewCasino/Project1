Din nya e-mailadress har blivit bekräftad och aktiverad.