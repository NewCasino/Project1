﻿Smart Underhållning
