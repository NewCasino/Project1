E-postadressen finns redan