﻿/game/gamerules.jsp?game=hrblackjackflash&lang=sv