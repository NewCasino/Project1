Ange ditt namn.