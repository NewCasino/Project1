Sofortbanking är ett lättanvändbart direktbetalningutförande med samma höga säkerhetsstandard som Internetbanken.