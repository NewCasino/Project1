﻿Fransk Roulette Serier
