﻿<!—Infoga Bakgrundsbild här -->
