Ditt efternamn innehåller otillåtna tecken