Neka