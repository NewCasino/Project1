﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Kasino Lobby
