Kontrollera att angivna uppgifter stämmer överens med uppgifterna för ditt AstroPay-kort.