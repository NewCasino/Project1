﻿Bonus ID


