Ange kontonumret.