﻿Abaqoos