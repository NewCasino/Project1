﻿Kort Nr.
