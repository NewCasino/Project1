Senaste vinnare: