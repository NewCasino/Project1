[Metadata:value(/Metadata/Settings.Operator_DisplayName)] Om oss