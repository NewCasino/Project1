Gratisspel