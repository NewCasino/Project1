﻿Nästa...

