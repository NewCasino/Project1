﻿
		The transaction could not be completed, may be due to connection problem. Click <a style="font-weight: bolder; text-decoration: none;" href="javascript:self.location.reload();">here</a> to retry.
        <br /><br />
        If the problem persist, please contact paysafecard <a style="font-weight: bolder; text-decoration: none;" href="http://www.paysafecard.com/uk/personal/contact-us/" target="_blank">support</a> or  go to <a style="font-weight: bolder; text-decoration: none;" href="https://customer.cc.at.paysafecard.com/psccustomer/GetWelcomePanelServlet?language=en" target="_blank">card’s balance page</a> to find out when the reserved amount will be available again.
	