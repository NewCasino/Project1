Stad/ort måste bestå av minst 2 tecken