﻿Mobilbetalning