Internt fel.