﻿Max.