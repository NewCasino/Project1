Kära  $USERNAME$, <br /><br />Detta e-postmeddelande får du för att bekräfta att ditt halvår av självutanförskapet har löpt ut och alla funktioner i ditt konto är nu aktiverat. <br /><br />Tveka inte att kontakta oss om ni har några frågor på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a><p> </p><p>Kind Hälsningar</p><p>[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Kund Support Teamet</p>