﻿/Metadata/Promotions
