﻿/game/gamerules.jsp?game=hrblackjack2-3h&lang=sv