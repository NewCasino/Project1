Uttag direkt till ditt NEOSURF konto