I menyn nedan kan du välja hur mycket du vill sätta in på ditt konto per dag, per vecka eller per månad. Dessa gränser är oberoende av gränserna eller de lägsta gränserna som erbjuds via metoderna på insättningssidan. När en gräns har angetts, får du ett bekräftelsemeddelande via e-post. Du kan minska din gräns när som helst via den här menyn. Men, om du vill ta bort eller öka din gräns tillämpas en väntetid på 7 dagar. Väntetiden ger dig tid att tänka över din ändring.