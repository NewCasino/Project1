Detta är ett automatiskt e-postmeddelande som du du kan svara på. <hr/><p>Kära $FIRSTNAME$</p><p>Ditt konto har spärrats på grund av alltför många ogiltiga inloggningsförsök och kommer automatiskt att öppnas upp igen efter 15 minuter..</p><p>Om du har glömt ditt lösenord och behöver ändra det, vänligen använd "Glömt lösenord"-länken på hemsidan.</p><p>för ytterligare hjälp kontakta<a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Vänliga Hälsningar, <br /> [Metadata:value(/Metadata/Settings.Operator_DisplayName)] Kundservice</p>