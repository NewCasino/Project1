﻿[Metadata:value(/Metadata/Settings.Operator_DisplayName)], Uteslutningslutningsperioden är över