Välj konto för debitering 