﻿Invalid user status