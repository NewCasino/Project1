﻿Kasino Lobby
