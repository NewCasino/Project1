Skriv