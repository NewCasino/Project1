﻿Totalt antal Casino FPP-poäng: 