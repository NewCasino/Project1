Spel som