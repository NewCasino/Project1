﻿[metadata:value(/TermsConditions/_Index_aspx.Title)]