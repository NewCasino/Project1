﻿Regler och villkor
