﻿Gräns:

