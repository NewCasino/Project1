Tack, din registrering är slutförd!