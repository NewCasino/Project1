﻿Yandex.Money
