Uttag av pengar direkt till ditt SOFORT-konto