Giropay är en betalningsmetod online som är fokuserad på den tyska marknaden. 