﻿<!—Infoga logga här -->
