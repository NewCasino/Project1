﻿Online chatt
