﻿<img src="//cdn.everymatrix.com/Shared/_files/Meddelande/få_mail_24x24.png" />
