Lägg till {0} i mina favoriter