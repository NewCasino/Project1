Mottagarens TC-nummer