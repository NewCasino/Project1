Ett år