﻿A technical error occurred. Invalid IP address. Please contact the merchant's customer service.