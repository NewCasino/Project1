AGMO är en ledande regional online-betaltjänstleverantör i CEE-regionen.