Den här transaktionen har avbrutits.