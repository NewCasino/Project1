Sydafrika, Rand