﻿EnterKontanter
