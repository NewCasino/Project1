Valideringskod