Online banköverföring