﻿<ol>
        
<li><strong>INTRODUKTION(UK License):</strong>
<p>
1.1.&nbsp;&nbsp; &nbsp; genom att använda och/eller besöka någon sektion av webbsidan [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] &nbsp; (the "Webbsidan"); eller öppna ett konto på webbsidan måste du acceptera:
<br/>
1.1.1.&nbsp;&nbsp; &nbsp;de allmäna villkoren, på den här sidan; 
<br/>
1.1.2.&nbsp;&nbsp; &nbsp;Integritetspolicy,
<br/>
1.1.3.&nbsp;&nbsp; &nbsp; alla spelregeler,
<br/>
1.1.4.&nbsp;&nbsp; &nbsp;alla villkor för&nbsp; kampanjer, bonusar och speciella erbjudanden kan hittas på webbsidan då och då.
<br/>
1.2.&nbsp;&nbsp; &nbsp;Alla villkoren ovanför ska tillsammans avses som "Villkoren".
<br/>
1.3.&nbsp;&nbsp; &nbsp;Varvänligen läs igenom villkoren noga innan du accepterar dem. Om du inte accepterar villkoren var snäll och öppna inte ett konto eller fortsätt på denna sida. Ditt fortsättande på denna sida accpeterar villkoren.
<br/>
1.4.&nbsp;&nbsp; &nbsp;Villkoren kommer att träda i kraft den 9:e Juni 2010.
</p>
</li>

<li><strong>PARTIES</strong>
<p>
2.1.&nbsp;&nbsp; &nbsp;Sportbok service och innehåll på den här webbsidan drivs av EveryMatrix Ltd, reg. no. C44411, 712, 14/19 Street, Valletta, VLT 1432 Malta. EveryMatrix underhåller och driver en fullständig hanterad Sportsbook, genom Letter of Intent Number LGA/CL2/497/2008 som utfärdats av the Maltese Lotteries och Gaming Authority under  Maltas lagar.
<br/>
2.2.&nbsp;&nbsp; &nbsp;References in Villkor om användning av  "oss", "vår," "vi" eller “Företaget” är refernser för den part som du har avtal med, som anges ovan.
</p>
</li>


<li><strong>ÄNDRING I VILLKORENS ANVÄNDNING</strong>
<p>
3.1.&nbsp;&nbsp; &nbsp;Vi kan behöva att ändra villkoren på grund av olika anledningar,även på grund av reklam, för att följa nya lagar eller regleringar i kundservices syfte. De nyaste villkoren kan nås här, och vilket datum de trädde i kraft.
<br/>
3.2.&nbsp;&nbsp; &nbsp;När vi gör ändringar i villkoren skulle vi vilja uppmärksamma dig om dessa, detta kommer vi att göra via e-post eller genom att lägga till en notis på webbsidan.
</p>
</li>


<li><strong>ÖPPNAR DITT KONTO</strong>
<p>
4.1.&nbsp;&nbsp; &nbsp;För att göra en satsning via webbsidan, måste du skapa ett konto på webbsidan ("Ditt Konto").
<br/>
4.2.&nbsp;&nbsp; &nbsp;på grund av olika juridiska och kommersiella skäl, tillåter vi inte att konton öppnas av eller används av kunder baserade eller domiclied i vissa jursidictions, inklusive USA. Om du är i en sådan jursidiction bör du inte skapa ett konto på denna webbsida eller använda den här webbsidan.
<br/>
4.3.&nbsp;&nbsp; &nbsp; För att öppna Ditt Konto för använding på den här webbsidan, kan du kontakta vår kundservice, eller genom att klicka <a href="/registrera">här</a> och följ instruktionerna på skärmen.
<br/>
4.4.&nbsp;&nbsp; &nbsp;När du öppnar Ditt Konto kommer duatt bli förfrågan att dela med dig av dina personligauppgifter, innefattar ditt namn, födelsedag, och lämpliga kontaktuppgifter, innefattade en adress, telefonnummer och e-postadress ("Dina Kontakuppgifter"). 
<br/>
4.5.&nbsp;&nbsp; &nbsp;Du är nu medvetenoch accepterar genom att använda webbsidans tillgångar att du kan både vinna och förlora pengar.
<br/>
4.6.&nbsp;&nbsp; &nbsp;Ditt Konto måste vara registreat som ditt eget, med korrekt namn. Du kan endast öppna ett konto för the sportsbook.Alla andra konton du skapar med oss relaterat till Servicen och webbsidan skall vara "Dubbla Konton" . Alla dubbel konton kan bli avstänga av oss direkt och:
<br/>
4.6.1.&nbsp;&nbsp; &nbsp;alla transaktioner utfördda från dubbel kontont kommer bli ogiltigt;
<br/>
4.6.2.&nbsp;&nbsp; &nbsp; Alla insater eller insätttningar gjorda på dubbel konton kommer lämnas tillbaka till dig; and
<br/>
4.6.3.&nbsp;&nbsp; &nbsp;eventuella vinster, eller bonusar som du har vunnit under tiden ditt dubbel konto var aktivt kommer att bli ogiltigt och kommer återlämnas till oss, och du måste lämna över alla pengar som har blivit uttagna från dubbel kontot
<br/>
4.7.&nbsp;&nbsp; &nbsp;Om du vill öppna ett annat konto, kan du kontatka Mangern på <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]" target="_blank">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>. Om ett nytt konto öppnas, stängs det gamla av.
<br/>
4.8.&nbsp;&nbsp; &nbsp;Du måste upprätthålla ditt konto och hålla personuppgifter uppdaterade.</p>
</li>


<li><strong>VERIFERING AV DIN INDENTIET;KRAVPÅ PENNINGTVÄTT</strong>
<p>
5.1.&nbsp;&nbsp; &nbsp;Garanterar du att:
<br/>
5.1.1.&nbsp;&nbsp; &nbsp;du inte är yngre än:
<br/>
5.1.1.1.&nbsp;&nbsp; &nbsp;18 (arton) år; or
<br/>
5.1.1.2.&nbsp;&nbsp; &nbsp;någon rättslig ålder vid spelande eller spelverksamhet enligt lag eller jurisdiktion som gäller kräver ("Laglig ålder"); att
<br/>
5.1.2.&nbsp;&nbsp; &nbsp;att dina uppgifter som du har lämnat in när du öppnar ditt konto är korrekt; och<br/>
5.1.3.&nbsp;&nbsp; &nbsp;Du är den rätta ägaren till ditt Konto.
<br/>
5.2.&nbsp;&nbsp; &nbsp;Genom att acceptera villkoren godkännr du även att vi gör olika verifierings undersökningar som vi kan behöva för oss själva eller om en tredje part behöver det (including, regulatory bodies) för att verifiera din intendiet och personuppgifter. ("Kontroller"). 
<br/>
5.3.&nbsp;&nbsp; &nbsp;Under tiden när vi gör kontroller så kan vi beränsa dina uttag från ditt spelkonto. 
<br/>
5.4.&nbsp;&nbsp; &nbsp;Under vissa omständigheter kan vi behöva kontakta dig för ytterligare information för att göra veriferingskontrollenfullständig. Om du inte kan ge oss ytterligare information så kan vi upphäva ditt konto eller göra en tillfällig avstängning till du har gett ytterligare information. Dessutom, måste du tillhandhålla identifikation varje gång du gör ett uttag värde av tvåtusentrehundra (EUR 2,300)eller.
<br/>
5.5.&nbsp;&nbsp; &nbsp;Om vi inte kan bekräfta att du inte över laglig ålder så kan vi stäng av Ditt Konto. Om det visar sig att du har spelat eller gjort några speltransaktioner,så:
<br/>
5.5.1.&nbsp;&nbsp; &nbsp;Kommer ditt Konto att bli avstängt;
<br/>
5.5.2.&nbsp;&nbsp; &nbsp;alla transaktioner du utförde undertidn du var minderårig kommer att ogiltighetförklaras, alla relaterade överföringar utfördart av dig kommer att bli återlämnat;
<br/>
5.5.3.&nbsp;&nbsp; &nbsp;alla satsningar för spel gjorda av dig under tiden du var minderårig kommer att lämnas tillbaka till dig; och<br/>
5.5.4.&nbsp;&nbsp; &nbsp;eventuella vinster som du har tillkommit under sådan tid kommer du att behöva betala böter för och du kommer att behöva lämna tillbaka alla uttag som har gjorts på ditt spelkonto till oss.</p>
</li>


<li><strong>ANVÄNDARNAMN, LÖSENORD, OCH KUNDINFORMATION</strong>
<p>
6.1.&nbsp;&nbsp; &nbsp;Efter att ha öppnat ett konto, är det inte tillåtet att överlämna (varken avsiktligt eller oavsiktligt) ditt användarnamn och lösenord till någon annan. Om du har förlorat eller glömt dina konto uppgifter kan du återfå ditt lösenord genom att klicka “Glömt lösenord” i länken under loggin portalen.</p>
</li>


<li><strong>INSÄTTNINGAR OCH UTTAG FRÅN DITT KONTO</strong>
<p>
7.1.&nbsp;&nbsp; &nbsp;Om du vill delta i någon satsningen eller spelande på webbsidan , måste du göra en insättning på ditt spelkonto som du kan använda för satsningar och spel. 
<br/>
7.2.&nbsp;&nbsp; &nbsp;Insättningar till och uttag från ett konto gjorda genom olika betalningsleverantörer kan ändrar då och då. Tillvägagångssätt, villkot och regler kan variera mellan olika betalningsleverantörer.Vi tar inte emot kontanter som skickas till oss. 
<br/>
7.3.&nbsp;&nbsp; &nbsp;Genom att överföra pengar tillåter du inte göra några återbetalningar eller upphänvande, om inte avsluta alla dina insättnigar in på ditt konto, och aceptera att göra en återbetalning till för obetalda insättningar.
<br/>
7.4.&nbsp;&nbsp; &nbsp;Ditt kontot är inte ett bankkonto, så därför har det ingen garanti, försäkran, sposerad eller skyddad av något banksystem. Insättningar hos oss på ditt konto kommer ha samma värde, alltså det kommer inte ske någon skillnad i värdet på din insättning. 
<br/>
7.5.&nbsp;&nbsp; &nbsp;Vi kan när som helst kvitta positiv balans på ditt konto mot eventuella belopp som du är skyldig oss när vi har startat om alla satsningar eller satsningar via dubbelkonto, maskopi, fusk, bedrägeri och kriminellverksamhet eller fel.
<br/>
7.6.&nbsp;&nbsp; &nbsp;Du är skyldig att rapportera dina vinster och förluster till ditt skatteverk och dina mydigheter.
<br/>
7.7.&nbsp;&nbsp; &nbsp;Du kan begära ett uttag av dina tillgångar från ditt konto när som helst under förutsättningen att:
<br/>
7.7.1.&nbsp;&nbsp; &nbsp;alla betalningar från ditt konto har blivit godkända och inget har blivit återkallat, eller avstängt;
<br/>
7.7.2.&nbsp;&nbsp; &nbsp;Alla kontroller som avses i punkt fem ovan har slutförts. 
<br/>
7.8.&nbsp;&nbsp; &nbsp;Alla godkända överföringar måste ha tillräcklig information, så som hur pengar ska bli överförda till dig.Vi kommer att hjälpa dig i dina frågor angående betalningsmetoder och valuta i dina överföringar. Detta, är dock inte garanetart. 
<br/>
7.9.&nbsp;&nbsp; &nbsp;Vi har rätten att ta en avgift enligt belopp för vår egna kostnader (inkluderat kosnaden vid överföringar) för uttag av pengar som inte har blivit insatta i något spel.
<br/>
7.10.1.Spelare som registerar sig med [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] måste göra en insättning från ett konto som är registrerat med dess egna namn.
<br/>
7.10.2.Vi tillåter inte tredje part insättningar, dvs, en vän, släkting, partner, make eller fru.
<br/>
7.10.3. Om vi upptäcker att detta har intäffat under våra rutin säkerhetskontroller, så kommer alla eventuella vinster att bli ogiltiga och kommer att skickas tillbaka till kasinot och ursprungs överföringen kommer att överföras till den rätte ägarens konto/bankkonto.
<br/>
7.10.5.Om överföring med masterkort inte är möjligt, måste kortinnehavaren fylla i ett 'kreditkorts verifering formulär' och skicka in identifikationsdokument till oss för att göra en verifiering.</p>
</li>


<li><strong>GÖRA EN SATSNING ELLER SPELA</strong>
<p>
8.1.&nbsp;&nbsp; &nbsp;Alla transtaktioner kommer att samlas på det språk som du valde för din trasaktion.
<br/>
8.2.&nbsp;&nbsp; &nbsp; Det är ditt ansvar att alla uppgifter för trasaktionerna är korrekta. 
<br/>
8.3.&nbsp;&nbsp; &nbsp;Du kan komma åt din transaktionshistorik på webbsidn.
<br/>
8.4.&nbsp;&nbsp; &nbsp;Vi har rätten att neka hela eller en del av dina transaktioner när som helst. Ingen transaktion är tillåten av oss, innan vi har bekräftat att du angett ett godkännande. Om du inte mottgit någon bekräftelse om att ni transaktion har blivit godkänd, bör du kontakta Kundsevice.
<br/>
8.5.&nbsp;&nbsp; &nbsp;När din satsning har blivit bekräftad, kan du inte avbryta transaktionen, utan vårt skriftliga medgivande.</p>
</li>


<li><strong>MASKOPI, FUSK, BEDRÄGERI OCH KRIMINELLVERKSAMHET</strong>
<p>
9.1.&nbsp;&nbsp; &nbsp;Följande handlingar är inte tillåtet och är en överträdle av villkoren:</p>
	<ul>
		<li>Maskopi med tredje part; </li>
		<li>ger en orättvis fördel eller påverkan (även känt som fusk), även utnutjanda av bedrägeri, kryphål eller fel i vår programvara använt automatiskt av spelare including the exploitation of a fault, loophole or error in our software, the use of automated players (ibland känd som 'robtspelare'); eller utnyttjande av ett 'fel';</li>
		<li>åtagande av bedrägerihandlingar för din fördel, även stulen, kopierad eller ogiltigt kredit- eller debitkort, som en finansieringskälla;</li>
		<li>Deltagande i något som helst kriminelverksamt, som pengatvätt och eller brott med kriminella konsekvenser.</li>
	</ul>
<p>
9.2.&nbsp;&nbsp; &nbsp;Vi tar ett ansvar för att förhindra sådana händelser; upptäcka dem och de relevanta spelarna;och ta itu med lämpliga valda spelare. Vi står inte för någon fölust eller skada som du eller någon annan spelare har ådrgit sig av maskopi, bedräger eller annan olagligverksamhet eller fusk, och annan handling kommer vi ha i vårt omdöme.
<br/>
9.3.&nbsp;&nbsp; &nbsp;Om du misstänker att en person utför maskopi, fusk eller bedrägeri, så bör du rappotera detta snarast genom att skicka ett e-post till oss.
<br/>
9.4.&nbsp;&nbsp; &nbsp;Vi har rätten att informera relevanta myndigeheter, andra spelbolag eller speloperatörer, andra serviceleverantörer och banker, kreditkortföretag,eletroniska betalningsleverantörer eller andra finasiella instutioner för din identier och för någon misstänk olaglig, bedrägare eller olämplig aktivit, och godkänner du att fullt ut samarbeta med oss att utreda sådana handlingar.</p>
</li>


<li><strong>ANDRA OTILLÅTNA HANDLINGAR</strong>
<p>
10.1.&nbsp;&nbsp; &nbsp;Du bör inte använda denna webbsida med ändamål är att kränka, missbruka, motbjuda,  rasistiskt, sexistiskt, diskriminera, eller stötande. Du får inte använda dig av ett kränkade eller aggrisivt språk eller biler; svordomar, hot, trakassera eller skällsord till någon annan, även andra spelare any other person, eller sådant beetende gentemot personalen på webbsidan och kundservicen.
<br/>
10.2.&nbsp;&nbsp; &nbsp; Du får inte korruptera webbsidan, flödet på webbsidan så det inte fungerar, eller använda dig av något som kan förhindra funktionen på webbsidan på något om helst vis, till exempel (men är inte begränsade) sprida virus, skapa oreda, "logic bombs" eller liknande. Flera svar eller "spam" är strikt förbjudet. Du får inte störa eller manipulera med, avlägsna eller på annat sätt ändra på något sätt någon information i någon form som ingår på webbplatsen.
<br/>
10.3.&nbsp;&nbsp; &nbsp;Du ska använda webbplatsen för personligt nöje och skall inte tillåtas att återskapa webbplatsen eller någon del av den i någon som helst form utan vårt medgivande.
<br/>
10.4.&nbsp;&nbsp; &nbsp;Du får inte försöka få obehörig åtkomst till webbplasten, serverna som lagars på webbsidan eller någon som helst server, dator eller databas ansluten till webbplatsen.Du får inte attackera webbplatsen genom en överbelastningsattack eller liknade. I händelse att bryta dessa bestämmelse kommer vi att anmäla detta brott till de relevanta brottbekämpande myndigheter och vi kommer att samarbeta med dessa myndigheter genom att avslöja din identiet till dem. I händelse av ett sådant brott, kommer din rätt att använda webbsidan omdelbart att upphöra.
<br/>
10.5.&nbsp;&nbsp; &nbsp;Vi tar inte något ansvar för någon förlut eller skada orsakad av en sprid överbelastningsattack, virus eller andra tekniskt skadliga matrial som kan ta skada på din datautrustning, datprogram, data eller andra materialpå grund av använding av webbsidan, din använding av webbplatsen eller nedladdnin av material som läggs på en sådan webbplats eller någon webbplats länkad till webbplatsen.
<br/>
10.6.&nbsp;&nbsp; &nbsp;Det ärförbjudet att sälja eller byta konton mellan spelare</p>
</li>


<li><strong>AVSTÄNGNING OCH UPPSÄGNING AV OSS</strong>
<p>
11.1.&nbsp;&nbsp; &nbsp;Det är företagspolicy i syfte av säkerheten och enligt sen maltesiska lagstifningen, att om ingen transaktion har registreats på ditt kono under trettio månder (ett “Inaktivt Konto”), Vi kommer att ge tillbaka saldot på kontot till dig. Om du inte kan lokalisera några tillgångarpå det kontot kommer det att överlämnas till Lotteries &amp; Gaming Authority of Malta. Alltså de tillgångar som finns tillgängliga för spelaren att ta utf.
<br/>
11.2.&nbsp;&nbsp; &nbsp;Ditt Inaktiva Konto kommer att bli avslutat i ett skriftligt meddelande (eller försök till meddelande) med hjälp av dina kontaktuppgifter. I händelse av en sådan uppsägning från oss, annat än om en sådan nedstäning och uppsägning görs i enlighet med punkt 11 (Maskopi, Fusk, Bedrägeri och kriminellverksamhet) eller punkt 20 (Brott mot användarvillkoren) med dessa villkor,kommer vi att betala tillbaka det saldo som finns på ditt konto. Om du inte kan lokaliseras, ska tillgångarna överföras till den berörda spelmyndigheten. </p>
</li>


<li><strong>ÄNDRING PÅ WEBBSIDAN</strong>
<p>
12.1.&nbsp;&nbsp; &nbsp;Vi kan i eget gottfinnande, ändra någon produkt som erbjuds via webbplatsen när som helst i syfte för att upprätthålla webbplatsen. &nbsp;</p>
</li>


<li><strong>IT FEL</strong>
<p>
13.1.&nbsp;&nbsp; &nbsp;När ett oväntat systemfel, fel eller fel som uppstår i software eller hårdvarasom vi använder för att tillhandahålla webbplatsen kommer vi att vidta omdelbara åtgärder för att lösa problemet. 
<br/>
13.2.&nbsp;&nbsp; &nbsp;Vi accepterar inte något IT-fel som orsakas av din utrustning som används för att få tillgång till webbplatsen eller som relaterar till din internetleverantör.</p>
</li>

<li><strong>FEL ELLER UTELÄMNINGAR</strong>
<p>
14.1.&nbsp;&nbsp; &nbsp;Ett antal omständigheter kan ett fel av oss uppstå när en satsning eller betalning görs. 
<br/>
14.2.&nbsp;&nbsp; &nbsp;[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)]  har rätten att avbryta en satsningen som är gjord på inkorrekta odds eller ombytta odds (där oddesen noteras mot fel lag) eller om satsningen är gjord efter ett event har startat och det är inte tillgängligt för livesatsningar. [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] har rätten att vägra, begränsa, stänga av eller sätta en grän på vilken satsnings som helst.
<br/>
14.3.&nbsp;&nbsp; &nbsp;Varken vi (inkluderat våra anställda och agenter) eller våra partners eller leverantörer ska vara ansvarig för eventuella förluster, inklusive förlut av vinster som är resultatet av något fel av oss eller fel av dig. Du kommer att förlora eventuella vinster/förluster som resulterar från sådan fel.</p>
</li>

<li><strong>UTESLUTNING PÅ VÅRT ANSVAR</strong>
<p>
15.1.&nbsp;&nbsp; &nbsp;Din tillång till användningen av produkter som erbjuds via webbplatsen är på egetbevåg och risk. 
<br/>
15.2.&nbsp;&nbsp; &nbsp;Vi kommer att förse webbsidan med rimliga färdigheter och omsorg och det väsentliga villkoren. We do not make any other promises or warranties the Website, or the products offered via the Website, and hereby exclude (to the extent permitted by law) all implied warranties in respect of the same.
<br/>
15.3.&nbsp;&nbsp; &nbsp;We shall not be liable to You in contract, tort (including negligence) or otherwise for any business losses, including but not limited to loss of data, profits, revenue, business, opportunity, goodwill, reputation or business interruption or for any losses which are not currently foreseeable by us arising out of the Terms of Use or Your use of the Website.</p>
</li>


<li><strong>BREACH OF THE TERMS OF USE</strong>
<p>
16.1.&nbsp;&nbsp; &nbsp; You shall compensate us in full for any claims, liabilities, costs, expenses (including legal fees) and any other charges that may arise as a result of your breach of the Terms.
<br/>
16.2.&nbsp;&nbsp; &nbsp;Where you are in material breach of the Terms, we reserve the right, but shall not be required, to:
<br/>
16.2.1.&nbsp;&nbsp; &nbsp;Provide you with notice (using Your Contact Details) that you are in breach requiring you to stop the relevant act or failure to act,
<br/>
16.2.2.&nbsp;&nbsp; &nbsp;suspend your Account so that you are unable to place bets or play games on the Website, 
<br/>
16.2.3.&nbsp;&nbsp; &nbsp; close Your Account with or without prior notice from us.
<br/>
16.2.4.&nbsp;&nbsp; &nbsp;recover from Your Account the amount of any pay-outs, bonuses or winnings which have been affected by any material breach.
<br/>
16.3.&nbsp;&nbsp; &nbsp;We have the right to disable any user identification code or password if in our reasonable opinion you have failed to comply with any of the provisions of the Terms.</p>
</li>


<li><strong>INTELLECTUAL PROPERTY RIGHTS</strong>
<p>
17.1.&nbsp;&nbsp; &nbsp;All website design, text, graphics, music, sound, photographs, video, the selection and arrangement thereof, software compilations, underlying source code, software and all other material contained within the Website are subject to copyright and other proprietary rights which are either owned by us or used under licence from third party rights owners. To the extent that any material contained on the Website may be downloaded or printed then such material may be downloaded to a single personal computer only and hard copy portions may be printed solely for your own personal and non-commercial use.
<br/>
17.2.&nbsp;&nbsp; &nbsp; Under no circumstances shall the use of the Website grant to any user any interest in any intellectual property rights (for example copyright, know-how or trade marks) owned by us or by any third party whatsoever.
<br/>
17.3.&nbsp;&nbsp; &nbsp;No rights whatsoever are granted to use or reproduce any trade names, trade marks or logos which appear on the Website except as specifically permitted in accordance with the Terms of Use.</p>
</li>


<li><strong>YOUR PERSONAL INFORMATION</strong>
<p>
18.1.&nbsp;&nbsp; &nbsp;We are required by law to comply with data protection requirements in the way in which we use any personal information collected from you in your use of the Website. We therefore take very seriously our obligations in relation to the way in which we use your personal information.
<br/>
18.2.&nbsp;&nbsp; &nbsp;By providing us with the information, you consent to our processing your personal Information for the purposes set out in the Term, for operating the Website or to comply with a legal or regulatory obligation.
<br/>
18.3.&nbsp;&nbsp; &nbsp;As a policy the Company will not disclose any personal information to anyone other than those employees that need access to your data to provide you with a service.
<br/>
18.4.&nbsp;&nbsp; &nbsp;We will retain copies of any communications that you send to us (including copies of any emails) in order to maintain accurate records of the information that we have received from you.</p>
</li>


<li><strong>USE OF COOKIES ON THE WEBSITE</strong>
<p>
19.1.&nbsp;&nbsp; &nbsp;The Website uses 'cookies' to assist the functionality of the Website. A cookie is a small file of text which is downloaded onto your computer when you access the Website and it allows us to recognise when you come back to the Website. Information on deleting or controlling cookies is available at www.aboutcookies.org. Please note that by deleting our cookies or disabling future cookies you may not be able to access certain areas or features of the Website.</p>
</li>


<li><strong>COMPLAINTS AND NOTICES</strong>
<p>
20.1.&nbsp;&nbsp; &nbsp;If You wish to make a complaint regarding the Website, a first step should be to, soon as reasonably possible, contact Customer Services.
<br/>
20.2.&nbsp;&nbsp; &nbsp;In the event of any dispute, you agree that the records of the server shall act as the final authority in determining the outcome of any claim.
<br/>
20.3.&nbsp;&nbsp; &nbsp;You agree that in the unlikely event of a disagreement between the result that appears on your screen and the game server, the result that appears on the game server will prevail, and you acknowledge and agree that our records will be the final authority in determining the terms and circumstances of your participation in the relevant online gaming activity and the results of this participation.
<br/>
20.4.&nbsp;&nbsp; &nbsp;When we wish to contact you regarding such a dispute, we will do so by using any of Your Contact Details.</p>
</li>


<li><strong>INTERPRETATION</strong>
<p>
21.1.&nbsp;&nbsp; &nbsp;The original text of the Terms is in English and any interpretation of them will be based on the original English text. If the Terms of Use or any documents or notices related to them are translated into any other language, the original English version will prevail.</p>
</li>


<li><strong>TRANSFER OF RIGHTS AND OBLIGATIONS</strong>
<p>
22.1.&nbsp;&nbsp; &nbsp;We reserve the right to transfer, assign, sublicense or pledge the Terms, in whole or in part, to any person, provided that any such assignment will be on the same terms or terms that are no less advantageous to You. </p>
</li>


<li><strong>EVENTS OUTSIDE OUR CONTROL</strong>
<p>
23.1.&nbsp;&nbsp; &nbsp; We will not be liable or responsible for any failure to perform, or delay in performance of, any of our obligations under the Terms of Use that is caused by events outside our reasonable control, including, without limitation, acts of God, war, civil commotion, interruption in public communications networks or services, industrial dispute or DDOS-attacks and similar Internet attacks having an adverse effect ("Force Majeure"). Our performance is deemed to be suspended for the period that the Force Majeure Event continues, and we will have an extension of time for performance for the duration of that period. We will use our reasonable endeavours to bring the Force Majeure Event to a close or to find a solution by which our obligations may be performed despite the Force Majeure Event.</p>
</li>


<li><strong>WAIVER</strong>
<p>
24.1.&nbsp;&nbsp; &nbsp;If we fail to insist upon strict performance of any of your obligations or if we fail to exercise any of the rights or remedies to which we are entitled, this shall not constitute a waiver of such rights or remedies and shall not relieve you from compliance with such obligations.
<br/>
24.2.&nbsp;&nbsp; &nbsp;A waiver by us of any default shall not constitute a waiver of any subsequent default. No waiver by us of any of the provisions of the Terms shall be effective unless it is expressly stated to be a waiver and is communicated to you in writing in accordance with above.</p>
</li>


<li><strong>SEVERABILITY</strong>
<p>
25.1.&nbsp;&nbsp; &nbsp;If any of the Terms are determined to be invalid, unlawful or unenforceable to any extent, such term, condition or provision will to that extent be severed from the remaining terms, conditions and provisions which will continue to be valid to the fullest extent permitted by law. In such cases, the part deemed invalid or unenforceable shall be amended in a manner consistent with the applicable law to reflect, as closely as possible, Our original intent.</p>
</li>


<li><strong>LAW AND JURISDICTION</strong>
<p>
26.1.&nbsp;&nbsp; &nbsp;The Terms of Use shall be governed by and interpreted in accordance with the laws of England and Wales save for any issues arising in respect to the Maltese licence which will be governed by Maltese Law in the Maltese Courts.
<br/>
26.2.&nbsp;&nbsp; &nbsp;The Courts of England and Wales shall have non-exclusive jurisdiction over any disputes arising out of the Terms of Use themselves.</p>
</li>


<li><strong>RESPONSIBLE GAMING AND GAMBLING</strong>
<p>
27.1.&nbsp;&nbsp; &nbsp;For those customers who wish to restrict their gambling, we provide a voluntary self-exclusion policy, which enables you to close Your Account or restrict your ability to place bets. If you require any information relating to this facility please speak to Customer Services.
<br/>
27.2.&nbsp;&nbsp; &nbsp;We will use our reasonable endeavours to ensure compliance with your self-exclusion. However you accept that we have no responsibility or liability whatsoever if you continue gambling and/or seek to use the Website and we fail to recognise or determine that.
<br/>
27.3.&nbsp;&nbsp; &nbsp;We are committed to supporting Responsible Gambling initiatives and encourage you to find information about Responsible Gambling at the websites of the following organisations:
<br/>
Gambling Therapy - www.gamblingtherapy.org
<br/>
Gordon House Association - 
<a href="http://www.gordonhouse.org.uk">www.gordonhouse.org.uk</a></p>
</li>

<li><strong>LINKS</strong>
<p>
28.1.&nbsp;&nbsp; &nbsp;Where we provide hyperlinks to other websites, we do so for information purposes only. You use any such links at your own risk and we accept no responsibility for the content or use of such websites, or for the information contained on them.</p>
</li>
    

</ol>

<p style="text-align:right">
    <button type="button" onclick="window.print(); return false" class="button button-print">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span>Print</span>
                </span>
            </span>
        </span>
    </button>
</p>

