Ange kontoinnehavarens filial.