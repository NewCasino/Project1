Ändra e-postadress