Om du är berättigad och har en bonuskod för bonus, ange koden nedan och klicka på "Skicka".