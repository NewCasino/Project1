Bank Transfer