﻿Det finns ett fel i din väns användarnamn eller E-post adress.
