Ogiltigt Ukash-värde.