Kortets utgivningsnummer