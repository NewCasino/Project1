Visa kreditkort