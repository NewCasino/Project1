<p>Hej $FIRSTNAME$,</p><p>Din utbetalning för $VOUCHERAMOUNT$ has been processed. har bearbetats. Nedan finns information om din kupong:</p><ul><li><strong>Ukash Kupong Nummer</strong>:$VOUCHERNUMBER$</li><li><strong>Ukash Kupong Summa</strong>:$VOUCHERAMOUNT$</li><li><strong>Ukash kupong förbrukningsdag </strong>:$VOUCHEREXPIRYDATE$</li></ul><p>Om du har några frågor angående din voucher vänligen tveka inte att kontakta <a href="mailto:[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]">[Metadata:htmlencode(/Metadata/Settings.Email_SupportAddress)]</a>.</p><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] teamet</p>