﻿Nedtrappning under 30 dagar
