Registrera ett nytt konto