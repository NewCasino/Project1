Postnummer