Ange ditt efternamn