Registrera ett Skrill-konto