Vänligen ange summa