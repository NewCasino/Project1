En 7-dagars uppehållsperiod, som bara kan användas två (2) gånger