Tonvis med sporthändelser pågår just nu!