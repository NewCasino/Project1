Betala per telefon (Tjekiska republiken)