Gör ett uttag direkt till ditt Yandex konto