﻿Antal Casino FPP poäng
