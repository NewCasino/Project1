﻿Casinospel - Teoretisk utbetalning