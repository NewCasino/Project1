Glömt lösenord