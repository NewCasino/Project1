Insättning {0} för {1} bonus!