Kortägarens namn behövs