﻿i-BANQ användar-MID krävs
