Det finns ingen aktiv bonus just nu