﻿Punto Banco Serier
