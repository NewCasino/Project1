 Fler bord 