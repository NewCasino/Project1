﻿Cool-off för 24 timmar
