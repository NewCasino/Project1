﻿Registreringen ej tillåten!
