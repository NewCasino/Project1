﻿/game/gamerules.jsp?game=lrblackjackpntn&lang=sv