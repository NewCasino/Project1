Kostnad