Från konto