Du kan inte göra uttag för att ditt konto inte är aktiverad