riktiga pengar