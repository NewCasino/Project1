﻿/game/gamerules.jsp?game=tribblemini&lang=sv