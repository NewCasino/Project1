Vänligen ange ditt namn