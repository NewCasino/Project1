﻿Nästa sida
