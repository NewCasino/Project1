Växlingsbelopp: