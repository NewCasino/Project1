Klicka för att visa kvittot för den här transaktionen.