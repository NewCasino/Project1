﻿Teoretisk vinståterbetalning
