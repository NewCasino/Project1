﻿Mata in ditt nya lösenord här
