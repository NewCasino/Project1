﻿/game/gamerules.jsp?game=txsholdem&lang=sv