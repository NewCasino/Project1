﻿Offline

