﻿felaktigt emailformat.
