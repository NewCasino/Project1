﻿Fel mobilnummer
