Mottagarens turkiska National ID