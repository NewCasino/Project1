Överför till bank