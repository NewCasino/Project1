Klicka för att visa spel från olika kategorier.