Lösenord