Landsprefix