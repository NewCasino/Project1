välj typ för din bonuskod