Betala per telefon (Italien)