Euro länder, Euro