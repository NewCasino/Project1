﻿Det tar bara 3 minuter
