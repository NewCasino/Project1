﻿Ditt efternamn måste innehålla minst 2 tecken
