Välj sorteringssätt...