Välj ditt riktnummer