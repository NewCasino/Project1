﻿Till
