﻿Konfiskera alla pengar på förverkade gods
