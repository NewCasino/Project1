Ogiltigt bankkontonummer