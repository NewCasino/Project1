﻿/game/gamerules.jsp?game=treypoker-1h&lang=sv