De nästkommande 3 månaderna