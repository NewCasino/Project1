﻿Vinnare
