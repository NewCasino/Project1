Ange ditt mobilnummer