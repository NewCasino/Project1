﻿Mobilprefix måste vara {0}.
