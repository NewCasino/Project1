﻿Casino Lobby
