﻿Spel Poäng
