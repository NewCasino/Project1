﻿Alltför många försök
