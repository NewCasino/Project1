Vänligen fyll i mottagarens TC nummer.