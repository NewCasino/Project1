﻿<style type="text/css">
.limit-overlay{display:none; position: fixed; top: 0; left: 0; z-index: 999998; background: #000; background:  rgba(0,0,0,0.8); filter: alpha(opacity=80);}
.limit-wrap{display:block; width:500px; height: 400px;color:#fff; background: #222; border:1px solid #999999; position: fixed; top: 200px; left: 0; z-index: 999999; }
.limit-box{display: block; margin: 40px auto; width: 70%;}
.limit-box h2{display: block; font-size: 24px; font-weight: bold; text-align: center; margin-bottom: 40px;}
.limit_item{display: block; font-size: 20px; line-height: 20px; margin: 20px 0; text-align: left;}
.limit_item label{margin-left: 20px;}
.limit-buttons{display: block; margin: 40px auto 0;}
</style>
