﻿Säkerhets svar
