Uttag direkt till ditt TELEINGRESO konto