﻿Live Multispelare Blackjack
