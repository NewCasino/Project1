Inkorrekt telefonnummer