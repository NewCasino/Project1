Gäller fr.o.m