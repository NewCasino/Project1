Inställning