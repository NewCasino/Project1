﻿Vilkor
