Skapa ett konto nu!