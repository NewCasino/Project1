﻿/game/gamerules.jsp?game=puntobanco&lang=sv