Tyvärr, du loggar in från ett land som vi inte accepterar insatser från. Vi kan inte slutföra din registrering.