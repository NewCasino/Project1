Captcha-koden är felaktig, försök igen.