﻿jackpot-spel
