Inte tillräckligt med pengar.