Beloppet överstiger den giltiga gränsen.