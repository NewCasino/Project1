Region/Stat