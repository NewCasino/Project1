﻿Gräns
