Filtrera spel efter tillverkare.