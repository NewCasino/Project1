﻿Classiska slots
