﻿Jag är missnöjd med sajten
