Du har avbrytit transaktionen