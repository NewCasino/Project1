Nästa {0} spel