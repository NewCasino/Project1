﻿Ta ut till ditt UIPAS-konto
