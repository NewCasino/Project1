﻿<ol>

    <li> <strong>Hur sätter jag in pengar på [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] Casino?</strong> 
        <p>
            Casino-saldot hålls separat från [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] huvudkontot så att du lätt får överblick, pengarna kan enkelt överföras mellan dessa två via funktionen "Överföring"&nbsp; som alltid visas på casinots högra sida när du är inloggad.
        </p>
    </li>

    <li> <strong>Hur rättvisa är spelen på er webbsida?</strong>
        <p>
            Vi försäkrar dig om att algoritmerna som används för att generera kort på vår webbsida är helt och hållet slumpmässiga. Våra spel är utvecklade med samma Sun Microsystem's Secure Random function för Java. Slumpgeneratorn och blandaren har utvecklats av en filosofie doktor inom matematik. Programvaran som vi använder för slumpmässiga spel har testats noggrant och har inte påvisat några metodfel eller förutsägbarhet, och har godkänts av eCOGRA.
        </p>
    </li>

    <li>
        <strong>Vad händer om ett spel blir avbrutet mitt i en spelrunda?</strong> 
        <p>
            Ställningen i varje spelrunda lagras automatiskt i systemets databas. Det säkerställer att ställningen i det senaste spelet som spelaren kunnat se alltid har lagrats och återupptas efter ett avbrott i systemet, internet eller serverfel, eller problem på kundens sida.
        </p>
    </li>

    <li>
        <strong>Hur många kortlekar finns det i Blackjack-spelet?</strong>
        <p>4 och 6 kortlekar används i våra Blackjack-spel.</p>
    </li>

    <li>
        <strong>Var hittar jag detaljerade anvisningar till era spel?</strong>
        <p>
            Alla våra spel har "Spelregler" på de specifika spelens egna sidor.
        </p>
    </li>

    <li>
        <strong>Hur mycket betalar webbsidan ut i genomsnitt?</strong>
        <p>
            Utbetalningarna varierar från spel till spel och över tid, men de teoretiska utbetalningarna ligger på cirka 97%. Utbetalningarna från spelen är hårdkodade och justeras inte av oss.
        </p>
    </li>

    <li>
        <strong>Kan jag prova spelen gratis?</strong>
        <p>
            Ja, du kan spela alla spel gratis om du väljer läget "Spela på skoj".
        </p>
    </li>

    <li>
        <strong>Kan jag ångar min insats efter att den&nbsp;  lagts på bordet?</strong>
        <p>
            Det kan vara möjligt innan spelet har startat men efter det att spelet har startat kan du inte ändra&nbsp; eller minska din insats.
        </p>
    </li>

    <li>
        <strong>Vad händer om min anslutning bryts under en spelrunda?</strong>
        <p>
            Spelet fortsätter från det läget det var i när du loggar in och öppnar spelet igen. Spelautomaterna som snurrade vid tiden för avbrottet slutförs även om anslutningen har brutits.
        </p>
    </li>

</ol>

<p style="text-align:right">
    <button type="button" onclick="window.print(); return false" class="button">
        <span class="button_Right">
            <span class="button_Left">
                <span class="button_Center">
                    <span>Print</span>
                </span>
            </span>
        </span>
    </button>
</p>