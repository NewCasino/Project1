﻿<p class="content"> Enligt våra licensregler satta av United Kingdom Gambling Commission (UKGC), [metadata:value(/Metadata/Settings.Operator_DisplayName)] måste vi informera dig att spelarmedel hålls på speciella 
Vid eventuell konkurs kommer spelarmedel anses tillhöra företagets tillgångar. Detta enligt UKGCs krav för segregering av konton som är separerade från företagets operativa konton.spelarmedel på basnivå. För mer info besök:</p>
     <a href="http://www.gamblingcommission.gov.uk/consumers/protection_of_customer_funds.aspx">www.gamblingcommission.gov.uk</a>

