﻿Jag har läst och godkänt den ovannämnda notifikationen
