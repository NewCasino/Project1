﻿Otillräckligt medel


