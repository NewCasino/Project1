Visa filtren för den här spellistan