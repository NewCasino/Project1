Transaktionen är inte slutförd, uppdatera den här sidan när transaktionen har slutförts.