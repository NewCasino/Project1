﻿eller

