Kompisens användarnamn