Visa den här guiden