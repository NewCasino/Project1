Problem med betalningar