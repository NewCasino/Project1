Spela med riktiga pengar