﻿Skräp
