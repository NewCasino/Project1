﻿/game/gamerules.jsp?game=fhvideopokerjob&lang=sv