Kontrollsiffra