﻿Tillbaka
