﻿US$ (USD)
