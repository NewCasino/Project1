﻿Virgin Islands(British)