Uttag direkt till ditt MULTIBANCO konto