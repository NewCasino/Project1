﻿/game/gamerules.jsp?game=hrscratchticketjp&lang=sv