﻿Ortfältet måste innehålla minst två tecken
