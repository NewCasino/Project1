﻿Välj din valuta
