Qiwi är en e-plånbok och terminalservice som erbjuder dig säkra betalningar online