﻿Your request could not be completed.Please call NETELLER (1-PAY) CustomerService at 86-13075600300 (nationwide mobile phone users), 86-108008530056(fixed line users - Northern China), 86-108001530056 (fixed line users - SouthernChina)