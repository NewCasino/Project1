﻿Steg 2. Överför <span style="font-weight: bold">{0}</span> <span style="font-weight: bold">{1}</span> till följande konto
