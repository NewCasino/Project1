Du får snart ett e-postmeddelande med ytterligare instruktioner för byte av lösenord.