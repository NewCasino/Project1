﻿Vänligen ange ditt namn
