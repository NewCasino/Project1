Fre