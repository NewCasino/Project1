﻿Affiliate kostnad