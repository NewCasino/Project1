Visa spel i alfabetisk ordning