﻿Överföringen lyckades.
