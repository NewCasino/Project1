Transaktionen har genomförts.