Kom ihåg 1 vecka