﻿Ort
