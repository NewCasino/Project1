Mitt favorit vad/bet?