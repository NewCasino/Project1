Ange ditt säkerhets-ID