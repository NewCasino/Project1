Lösenordet får inte vara samma som användarnamnet