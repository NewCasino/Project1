Visa favoritbord