﻿CreditMisslyckades