﻿Falsk
