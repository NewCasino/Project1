<p>När pengarna mottagits och godkänts kommer vi kreditera ditt spelkonto. Du behöver då följande detaljer när du ska göra en banköverföring </p><p>Vänligen gör betalning till  <ul> <li> <strong>Kontoägare</strong> : OddsMatrix Ltd</li> <li> <strong>Ägares adress</strong> : Vincenti Buildings, Suite 713, 14/19 Strait Street, Valletta, VLT 1432, Malta</li> <li> <strong>Bank name</strong> : Bank of Valletta</li> <li> <strong>Bank address</strong> : 86, South Street, Valletta VLT 1105-Malta</li> <li> <strong>SWIFT</strong> : VALLMTMT</li> </ul></p> <p>Below are IBAN numbers for each currency<ul><li> <strong>EUR</strong> MT25VALL22013000000040018502408</li><li> <strong>SEK</strong> MT11VALL22013000000040018502466</li><li> <strong>DKK</strong> MT34VALL22013000000040018502440</li><li> <strong>USD</strong> MT04VALL22013000000040018502495</li><li> <strong>GBP</strong> MT73VALL22013000000040018510759</li><li> <strong>NOK</strong> MT73VALL22013000000040018502453</li><li> <strong>PLN</strong> MT73VALL22013000000040019112062</li><li> <strong>CZK</strong> MT13VALL22013000000040019112075</li></ul></p><p> Vänligen notera att vi inte kommer att debitera dig för att du använder banköverföring, men vi rekommenderar dig att kontollera med din bank om de har några avgifter som de kan debitera dig för. </p>