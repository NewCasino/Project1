﻿Huvudmeny
