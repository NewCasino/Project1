﻿/game/gamerules.jsp?game=roulette2adv&lang=sv