Börja satsa på sporter 