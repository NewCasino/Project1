﻿Bonuskod
