﻿Dina inställningar har sparats
