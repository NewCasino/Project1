﻿<!—Infoga Logga här -->
