﻿Ukash-nummer