Det bekräftande e-mailet har skickats till din nya e-post inkorg, vänligen titta i din inkorg och aktivera den nya e-postadressen.