Clearingnummer