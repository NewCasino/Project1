Under 18 år