﻿Byt lösenord