Uttag av pengar direkt till ditt ABAQOOS-konto