﻿Toggle

