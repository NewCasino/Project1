﻿Referens
