Uttag av pengar direkt till ditt TrustPay-konto