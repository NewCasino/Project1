arabiska