﻿klassiset-kolikkopelit
