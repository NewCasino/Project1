Dealerns namn