﻿Skriv

