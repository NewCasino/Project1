Betalning via mobil