I kö