﻿Bankkonto
