Fel, det här spelet är inte tillgängligt längre!