﻿/game/gamerules.jsp?game=zodiac&lang=sv