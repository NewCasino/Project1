Uttag pågår