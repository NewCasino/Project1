Behandlar debitering