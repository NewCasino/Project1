Helskärm