﻿Neteller(Grekland)
