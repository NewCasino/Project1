Varianter: