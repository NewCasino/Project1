﻿Blackjack Serier
