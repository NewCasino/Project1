﻿Spela och gå
