Om du vill begränsa ditt spelande och göra ett uppehåll, ger vi dig följande möjligheter:<br>
Spärra min inloggning under