Filialkod