Uttag av pengar direkt till ditt Moneta-konto