﻿/game/gamerules.jsp?game=crusaders&lang=sv