Välj ett bankkonto