Du måste vara över {0} år