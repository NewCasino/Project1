Visa Debet