﻿Din mobil stöds inte av den valda banken, vänligen uppdatera din mobil för att fortsätta med insättningen

