﻿Deposit To