﻿Mikrospelning
