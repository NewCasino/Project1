﻿Andra spel
