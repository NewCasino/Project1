<p>Hej $FIRSTNAME$,</p><p>Tack för att du kontaktar [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)], Vi har tagit emot din begäran gällande ditt bortglömda lösenord. Klicka på följande länk för att återställa ditt lösenord. </p><p><a href="$RESETLINK$">$RESETLINK$</a></p><p>Denna länk är giltig i 24 timmar och kan bara användas en gång<p><p>Om du inte vill ändra ditt lösenord kan du ignorera detta mail <p/><p>Hälsningar,<br /> [Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] team</p>