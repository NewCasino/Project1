﻿Svenska kronor (SEK)
