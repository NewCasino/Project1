Skriv in tecknen på bilden.