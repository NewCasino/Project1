﻿Meddelandet har sänts. Vi kommer att återkomma till dig så snart som möjligt.

