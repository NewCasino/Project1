﻿BOCASH-kod