Om du har frågor, klicka här för att kontakta kundtjänst.