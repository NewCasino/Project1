﻿Credit Card
