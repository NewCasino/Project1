﻿/game/gamerules.jsp?game=blackjackmini&lang=sv