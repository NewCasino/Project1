Ett 1 års självutslutningsperiod