Gör ett uttag direkt med ditt Georgian Card