﻿Öppna Konto
