Uttag av pengar direkt till ditt PAGOFACIL-konto