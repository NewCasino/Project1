Uttag direkt till ditt Voucher konto