﻿/game/gamerules.jsp?game=jacksorbetter50&lang=sv