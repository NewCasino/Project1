﻿Otillgänglig bank
