Ange bordets namn: