Du kan för tillfället inte ändra din e-mail adress då ditt konto är inaktiverat. Ett e-mail för att aktivera ditt konto har skickats till den e-mailadress du använde vid registrering. Vänligen klicka på länken i e-mailet för att aktivera ditt konto. Om du inte får e-mailet var vänlig kontakta <a href="mailto:[Metadata:value(/Metadata/Settings.Email_SupportAddress)]">[Metadata:value(/Metadata/Settings.Email_SupportAddress)]</a>.