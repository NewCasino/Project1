﻿Användarnamnet redan upptaget
