﻿/game/gamerules.jsp?game=vault&lang=sv