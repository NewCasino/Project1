﻿Mottagarens namn
