Det är ett säkert och bekvämt sätt att spendera pengar online.