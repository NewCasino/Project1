Hitta en kompis via användarnamn.