﻿Bonus summa