Din kompis konto är blockerat.