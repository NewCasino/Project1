Väntande uttag