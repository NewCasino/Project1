﻿Skicka verifieringskod

