﻿Neteller(Austria)