Meddelandet har skickats och vi återkommer till dig så snart som möjligt.