[Metadata:htmlencode(/Metadata/Settings.Operator_DisplayName)] -Bekräftning på ändring av e-mailadress