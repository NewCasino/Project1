﻿/game/gamerules.jsp?game=lrtreypoker-1h&lang=sv