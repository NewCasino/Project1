Ogiltigt e-post format