Länken är felaktig eller har löpt ut.