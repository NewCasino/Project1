﻿POLi