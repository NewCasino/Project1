﻿Kreditkort
